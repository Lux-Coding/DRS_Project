--------------------------------------------------------------------------------
-- Title       : Write parallel digital audio data stream into a .wav file
-- Project     : FPGA Based Digital Signal Processing
--               FH OÖ Hagenberg/HSD, SCD5
--------------------------------------------------------------------------------
-- RevCtrl     : $Id: ParToWav-e.vhd 704 2017-10-27 19:25:59Z mroland $
-- Authors     : Markus Pfaff, Linz/Austria, Copyright (c) 2003-2005
--               Michael Roland, Hagenberg/Austria, Copyright (c) 2011-2017
--------------------------------------------------------------------------------
-- Description : Not intended for synthesis!
--               After the input wave is at its end the unit will write
--               additional samples into the WavOutFile. This is only done with
--               valid samples (i.e. the valid line has to be activated to flag
--               the sample valid).
--               
--               A problem with writing a .wav file: when writing a .wav file
--               the length of the file must be known from the beginning,
--               because the chunks contain their own lengths as explicit values
--               right at the start of the chunk. Thus the whole file content
--               has to be known before writing the file.
--               
--               Solution: A raw file is written simultaneously with simulation
--               progress. Under the circumstances stated below this raw file is
--               converted into a valid .wav file.
--               
--               Two questions arise:
--               - When simulating through a whole input .wav file: When is it
--                 at its end?
--                 Solution: The .wav file player (A/D converter model) has to
--                 signal the end of its input file to the sample receiver (D/A
--                 converter model).
--               - After the wave input to the DSP has ended the output of the
--                 DSP might still be of interest for some further time. For
--                 example when a delay algorithm is implemented the delay will
--                 last longer than the input wave. The wave file written to
--                 disk should therefore keep on for some extra time.
--               - When the user wants to hear the sound before the simulation
--                 is at its end: how to manage versions in between that are
--                 valid .wav files?
--                 Solution: Force the signal that flags the end of the input
--                 .wav file to its active value. The model will then convert
--                 the raw file as it is up to now in a valid .wav file.
--                 Afterwards the model suspends forever, i.e. the .wav file
--                 cannot be written a second time.
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.Global.all;
use work.RiffFileTreatment.all;

entity ParToWav is
  
  generic (
    gWavFileName                 : string := "./WetResult.wav";
    gRawWavFileName              : string := "./WetRawResult.raw";
    -- After the wave has ended it might be interesting to record the
    -- output of the DSP section for some further time. This will be
    -- especially interesting if the DSP section delays the signal.
    gRecordingDurationAftWaveEnd : time   := 2 ms;
    -- Parameters for .wav file. These parameters are taken by the model
    -- as-is and written into the created .wav file without modification.
    -- Thus, a reader of the .wav file generated by this model will always
    -- trust that the data found in the file matches these parameters
    -- (even if it doesn't). The user of the model has to assure that the
    -- parameters are adjusted correctly.
    gFormatTag                   : aWord  := 1;
    -- Word length of audio data at the interface
    gAudioBitWidth               : aWord  := cDefaultAudioBitWidth;
    -- Word length of audio data in the .wav file
    gWavFileBitWidth             : aWord  := 16;
    gChannels                    : aWord  := 2;
    gSampleRate                  : aDword := 44100); -- in Hz

  port (
    iClk : in std_ulogic;

    iDL, iDR     : in aAudioData(0 downto -(gAudioBitWidth-1));
    iValL, iValR : in std_ulogic;

    -- Controlling the model: Conversion of the .raw
    -- file into the .wav file is started when this input transits from
    -- false to true.
    iWaveAtEnd : in boolean := false);

begin

  assert gFormatTag = 1
    report "Mp: Only WAVE format 1 (Microsoft PCM) can be written."
    severity failure;

  assert gChannels = 2
    report "Mp: Only stereo .wav files can be written."
    severity failure;

  assert gWavFileBitWidth = 16
    report "Mp: Only audio data of 16 bit word length can be written."
    severity failure;

  assert (gSampleRate = 44100)
    or (gSampleRate = 48000)
    or (gSampleRate = 88200)
    or (gSampleRate = 96000)
    report "Mp: Using the non standard sample rate of " & aDword'image(gSampleRate) & " Hz."
    severity warning;

end ParToWav;

