-- Copyright (C) 2018  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details.

-- VENDOR "Altera"
-- PROGRAM "Quartus Prime"
-- VERSION "Version 18.1.0 Build 625 09/12/2018 SJ Lite Edition"

-- DATE "12/12/2021 02:42:30"

-- 
-- Device: Altera 5CSEMA5F31C6 Package FBGA896
-- 

-- 
-- This VHDL file should be used for ModelSim (VHDL) only
-- 

LIBRARY ALTERA;
LIBRARY ALTERA_LNSIM;
LIBRARY CYCLONEV;
LIBRARY IEEE;
USE ALTERA.ALTERA_PRIMITIVES_COMPONENTS.ALL;
USE ALTERA_LNSIM.ALTERA_LNSIM_COMPONENTS.ALL;
USE CYCLONEV.CYCLONEV_COMPONENTS.ALL;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY 	TbdRxFskBasic IS
    PORT (
	iClk : IN std_logic;
	inResetAsync : IN std_logic;
	iSwitch : IN IEEE.STD_LOGIC_1164.std_ulogic_vector(9 DOWNTO 0);
	inButton : IN IEEE.STD_LOGIC_1164.std_ulogic_vector(3 DOWNTO 1);
	oSEG0 : OUT IEEE.STD_LOGIC_1164.std_ulogic_vector(6 DOWNTO 0);
	oSEG1 : OUT IEEE.STD_LOGIC_1164.std_ulogic_vector(6 DOWNTO 0);
	oSEG2 : OUT IEEE.STD_LOGIC_1164.std_ulogic_vector(6 DOWNTO 0);
	oSEG3 : OUT IEEE.STD_LOGIC_1164.std_ulogic_vector(6 DOWNTO 0);
	oSEG4 : OUT IEEE.STD_LOGIC_1164.std_ulogic_vector(6 DOWNTO 0);
	oSEG5 : OUT IEEE.STD_LOGIC_1164.std_ulogic_vector(6 DOWNTO 0);
	oLed : OUT IEEE.STD_LOGIC_1164.std_ulogic_vector(9 DOWNTO 0);
	oI2cSclk : OUT std_logic;
	ioI2cSdin : INOUT std_logic;
	oMclk : OUT std_logic;
	oBclk : OUT std_logic;
	iADCdat : IN std_logic;
	oDACdat : OUT std_logic;
	oADClrc : OUT std_logic;
	oDAClrc : OUT std_logic
	);
END TbdRxFskBasic;

-- Design Ports Information
-- iSwitch[1]	=>  Location: PIN_AC12,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: Default
-- iSwitch[2]	=>  Location: PIN_AF9,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: Default
-- iSwitch[3]	=>  Location: PIN_AF10,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: Default
-- iSwitch[4]	=>  Location: PIN_AD11,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: Default
-- iSwitch[5]	=>  Location: PIN_AD12,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: Default
-- iSwitch[6]	=>  Location: PIN_AE11,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: Default
-- iSwitch[7]	=>  Location: PIN_AC9,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: Default
-- iSwitch[8]	=>  Location: PIN_AD10,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: Default
-- iSwitch[9]	=>  Location: PIN_AE12,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: Default
-- inButton[1]	=>  Location: PIN_AA15,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: Default
-- inButton[2]	=>  Location: PIN_W15,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: Default
-- inButton[3]	=>  Location: PIN_Y16,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: Default
-- oSEG0[0]	=>  Location: PIN_AE26,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oSEG0[1]	=>  Location: PIN_AE27,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oSEG0[2]	=>  Location: PIN_AE28,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oSEG0[3]	=>  Location: PIN_AG27,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oSEG0[4]	=>  Location: PIN_AF28,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oSEG0[5]	=>  Location: PIN_AG28,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oSEG0[6]	=>  Location: PIN_AH28,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oSEG1[0]	=>  Location: PIN_AJ29,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oSEG1[1]	=>  Location: PIN_AH29,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oSEG1[2]	=>  Location: PIN_AH30,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oSEG1[3]	=>  Location: PIN_AG30,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oSEG1[4]	=>  Location: PIN_AF29,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oSEG1[5]	=>  Location: PIN_AF30,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oSEG1[6]	=>  Location: PIN_AD27,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oSEG2[0]	=>  Location: PIN_AB23,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oSEG2[1]	=>  Location: PIN_AE29,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oSEG2[2]	=>  Location: PIN_AD29,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oSEG2[3]	=>  Location: PIN_AC28,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oSEG2[4]	=>  Location: PIN_AD30,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oSEG2[5]	=>  Location: PIN_AC29,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oSEG2[6]	=>  Location: PIN_AC30,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oSEG3[0]	=>  Location: PIN_AD26,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oSEG3[1]	=>  Location: PIN_AC27,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oSEG3[2]	=>  Location: PIN_AD25,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oSEG3[3]	=>  Location: PIN_AC25,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oSEG3[4]	=>  Location: PIN_AB28,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oSEG3[5]	=>  Location: PIN_AB25,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oSEG3[6]	=>  Location: PIN_AB22,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oSEG4[0]	=>  Location: PIN_AA24,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oSEG4[1]	=>  Location: PIN_Y23,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oSEG4[2]	=>  Location: PIN_Y24,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oSEG4[3]	=>  Location: PIN_W22,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oSEG4[4]	=>  Location: PIN_W24,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oSEG4[5]	=>  Location: PIN_V23,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oSEG4[6]	=>  Location: PIN_W25,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oSEG5[0]	=>  Location: PIN_V25,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oSEG5[1]	=>  Location: PIN_AA28,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oSEG5[2]	=>  Location: PIN_Y27,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oSEG5[3]	=>  Location: PIN_AB27,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oSEG5[4]	=>  Location: PIN_AB26,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oSEG5[5]	=>  Location: PIN_AA26,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oSEG5[6]	=>  Location: PIN_AA25,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oLed[0]	=>  Location: PIN_V16,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oLed[1]	=>  Location: PIN_W16,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oLed[2]	=>  Location: PIN_V17,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oLed[3]	=>  Location: PIN_V18,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oLed[4]	=>  Location: PIN_W17,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oLed[5]	=>  Location: PIN_W19,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oLed[6]	=>  Location: PIN_Y19,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oLed[7]	=>  Location: PIN_W20,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oLed[8]	=>  Location: PIN_W21,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oLed[9]	=>  Location: PIN_Y21,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oI2cSclk	=>  Location: PIN_J12,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oMclk	=>  Location: PIN_G7,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oBclk	=>  Location: PIN_H7,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oDACdat	=>  Location: PIN_J7,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oADClrc	=>  Location: PIN_K8,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- oDAClrc	=>  Location: PIN_H8,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- ioI2cSdin	=>  Location: PIN_K12,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: 16mA
-- iClk	=>  Location: PIN_AF14,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: Default
-- inResetAsync	=>  Location: PIN_AA14,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: Default
-- iSwitch[0]	=>  Location: PIN_AB12,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: Default
-- iADCdat	=>  Location: PIN_K7,	 I/O Standard: 3.3-V LVTTL,	 Current Strength: Default


ARCHITECTURE structure OF TbdRxFskBasic IS
SIGNAL gnd : std_logic := '0';
SIGNAL vcc : std_logic := '1';
SIGNAL unknown : std_logic := 'X';
SIGNAL devoe : std_logic := '1';
SIGNAL devclrn : std_logic := '1';
SIGNAL devpor : std_logic := '1';
SIGNAL ww_devoe : std_logic;
SIGNAL ww_devclrn : std_logic;
SIGNAL ww_devpor : std_logic;
SIGNAL ww_iClk : std_logic;
SIGNAL ww_inResetAsync : std_logic;
SIGNAL ww_iSwitch : std_logic_vector(9 DOWNTO 0);
SIGNAL ww_inButton : std_logic_vector(3 DOWNTO 1);
SIGNAL ww_oSEG0 : std_logic_vector(6 DOWNTO 0);
SIGNAL ww_oSEG1 : std_logic_vector(6 DOWNTO 0);
SIGNAL ww_oSEG2 : std_logic_vector(6 DOWNTO 0);
SIGNAL ww_oSEG3 : std_logic_vector(6 DOWNTO 0);
SIGNAL ww_oSEG4 : std_logic_vector(6 DOWNTO 0);
SIGNAL ww_oSEG5 : std_logic_vector(6 DOWNTO 0);
SIGNAL ww_oLed : std_logic_vector(9 DOWNTO 0);
SIGNAL ww_oI2cSclk : std_logic;
SIGNAL ww_oMclk : std_logic;
SIGNAL ww_oBclk : std_logic;
SIGNAL ww_iADCdat : std_logic;
SIGNAL ww_oDACdat : std_logic;
SIGNAL ww_oADClrc : std_logic;
SIGNAL ww_oDAClrc : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~8_ACLR_bus\ : std_logic_vector(1 DOWNTO 0);
SIGNAL \TheRxFsk|Lowpass|Mult0~8_CLK_bus\ : std_logic_vector(2 DOWNTO 0);
SIGNAL \TheRxFsk|Lowpass|Mult0~8_ENA_bus\ : std_logic_vector(2 DOWNTO 0);
SIGNAL \TheRxFsk|Lowpass|Mult0~8_AX_bus\ : std_logic_vector(17 DOWNTO 0);
SIGNAL \TheRxFsk|Lowpass|Mult0~8_AY_bus\ : std_logic_vector(18 DOWNTO 0);
SIGNAL \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\ : std_logic_vector(63 DOWNTO 0);
SIGNAL \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTADATAIN_bus\ : std_logic_vector(39 DOWNTO 0);
SIGNAL \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTAADDR_bus\ : std_logic_vector(6 DOWNTO 0);
SIGNAL \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBADDR_bus\ : std_logic_vector(6 DOWNTO 0);
SIGNAL \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\ : std_logic_vector(39 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_AX_bus\ : std_logic_vector(17 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_AY_bus\ : std_logic_vector(18 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\ : std_logic_vector(63 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_AX_bus\ : std_logic_vector(17 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_AY_bus\ : std_logic_vector(18 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\ : std_logic_vector(63 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_AX_bus\ : std_logic_vector(17 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_AY_bus\ : std_logic_vector(18 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\ : std_logic_vector(63 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_AX_bus\ : std_logic_vector(17 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_AY_bus\ : std_logic_vector(18 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\ : std_logic_vector(63 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a0_PORTAADDR_bus\ : std_logic_vector(8 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a0_PORTADATAOUT_bus\ : std_logic_vector(19 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a4_PORTAADDR_bus\ : std_logic_vector(8 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a4_PORTADATAOUT_bus\ : std_logic_vector(19 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTADATAIN_bus\ : std_logic_vector(19 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTAADDR_bus\ : std_logic_vector(8 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBADDR_bus\ : std_logic_vector(8 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\ : std_logic_vector(19 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a4_PORTADATAIN_bus\ : std_logic_vector(19 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a4_PORTAADDR_bus\ : std_logic_vector(8 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a4_PORTBADDR_bus\ : std_logic_vector(8 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a4_PORTBDATAOUT_bus\ : std_logic_vector(19 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a0_PORTAADDR_bus\ : std_logic_vector(8 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a0_PORTADATAOUT_bus\ : std_logic_vector(19 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a12_PORTAADDR_bus\ : std_logic_vector(8 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a12_PORTADATAOUT_bus\ : std_logic_vector(19 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTADATAIN_bus\ : std_logic_vector(19 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTAADDR_bus\ : std_logic_vector(8 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBADDR_bus\ : std_logic_vector(8 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\ : std_logic_vector(19 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a12_PORTADATAIN_bus\ : std_logic_vector(19 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a12_PORTAADDR_bus\ : std_logic_vector(8 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a12_PORTBADDR_bus\ : std_logic_vector(8 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a12_PORTBDATAOUT_bus\ : std_logic_vector(19 DOWNTO 0);
SIGNAL \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_VCOPH_bus\ : std_logic_vector(7 DOWNTO 0);
SIGNAL \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_MHI_bus\ : std_logic_vector(7 DOWNTO 0);
SIGNAL \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~PLL_REFCLK_SELECT_CLKIN_bus\ : std_logic_vector(3 DOWNTO 0);
SIGNAL \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~PLL_RECONFIG_MHI_bus\ : std_logic_vector(7 DOWNTO 0);
SIGNAL \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~PLL_RECONFIG_SHIFTEN_bus\ : std_logic_vector(8 DOWNTO 0);
SIGNAL \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~PLL_OUTPUT_COUNTER_VCO0PH_bus\ : std_logic_vector(7 DOWNTO 0);
SIGNAL \TheRxFsk|Lowpass|Mult0~40\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~41\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~42\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~43\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~44\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~45\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~46\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~47\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~48\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~49\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~50\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~51\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~52\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~53\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~54\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~55\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~56\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~57\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~58\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~59\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~60\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~61\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~62\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~63\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~64\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~65\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~66\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~67\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~68\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~69\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~70\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~71\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~40\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~41\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~42\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~43\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~44\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~45\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~46\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~47\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~48\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~49\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~50\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~51\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~52\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~53\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~54\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~55\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~56\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~57\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~58\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~59\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~60\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~61\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~62\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~63\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~64\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~65\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~66\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~67\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~68\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~69\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~70\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~71\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~40\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~41\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~42\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~43\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~44\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~45\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~46\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~47\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~48\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~49\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~50\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~51\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~52\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~53\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~54\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~55\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~56\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~57\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~58\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~59\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~60\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~61\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~62\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~63\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~64\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~65\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~66\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~67\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~68\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~69\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~70\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~71\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~40\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~41\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~42\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~43\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~44\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~45\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~46\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~47\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~48\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~49\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~50\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~51\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~52\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~53\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~54\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~55\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~56\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~57\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~58\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~59\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~60\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~61\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~62\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~63\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~64\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~65\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~66\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~67\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~68\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~69\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~70\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~71\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~40\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~41\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~42\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~43\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~44\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~45\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~46\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~47\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~48\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~49\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~50\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~51\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~52\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~53\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~54\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~55\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~56\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~57\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~58\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~59\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~60\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~61\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~62\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~63\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~64\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~65\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~66\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~67\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~68\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~69\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~70\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~71\ : std_logic;
SIGNAL \iSwitch[1]~input_o\ : std_logic;
SIGNAL \iSwitch[2]~input_o\ : std_logic;
SIGNAL \iSwitch[3]~input_o\ : std_logic;
SIGNAL \iSwitch[4]~input_o\ : std_logic;
SIGNAL \iSwitch[5]~input_o\ : std_logic;
SIGNAL \iSwitch[6]~input_o\ : std_logic;
SIGNAL \iSwitch[7]~input_o\ : std_logic;
SIGNAL \iSwitch[8]~input_o\ : std_logic;
SIGNAL \iSwitch[9]~input_o\ : std_logic;
SIGNAL \inButton[1]~input_o\ : std_logic;
SIGNAL \inButton[2]~input_o\ : std_logic;
SIGNAL \inButton[3]~input_o\ : std_logic;
SIGNAL \~QUARTUS_CREATED_GND~I_combout\ : std_logic;
SIGNAL \iClk~input_o\ : std_logic;
SIGNAL \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~PLL_REFCLK_SELECT_O_EXTSWITCHBUF\ : std_logic;
SIGNAL \inResetAsync~input_o\ : std_logic;
SIGNAL \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~PLL_REFCLK_SELECT_O_CLKOUT\ : std_logic;
SIGNAL \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_MHI2\ : std_logic;
SIGNAL \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_MHI3\ : std_logic;
SIGNAL \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_MHI4\ : std_logic;
SIGNAL \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_MHI5\ : std_logic;
SIGNAL \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_MHI6\ : std_logic;
SIGNAL \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_MHI7\ : std_logic;
SIGNAL \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~PLL_RECONFIG_O_UP\ : std_logic;
SIGNAL \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_MHI1\ : std_logic;
SIGNAL \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~PLL_RECONFIG_O_SHIFTENM\ : std_logic;
SIGNAL \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_MHI0\ : std_logic;
SIGNAL \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~PLL_RECONFIG_O_SHIFT\ : std_logic;
SIGNAL \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_CNTNEN\ : std_logic;
SIGNAL \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~PLL_RECONFIGSHIFTEN6\ : std_logic;
SIGNAL \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_TCLK\ : std_logic;
SIGNAL \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_VCOPH0\ : std_logic;
SIGNAL \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_VCOPH1\ : std_logic;
SIGNAL \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_VCOPH2\ : std_logic;
SIGNAL \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_VCOPH3\ : std_logic;
SIGNAL \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_VCOPH4\ : std_logic;
SIGNAL \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_VCOPH5\ : std_logic;
SIGNAL \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_VCOPH6\ : std_logic;
SIGNAL \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_VCOPH7\ : std_logic;
SIGNAL \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\ : std_logic;
SIGNAL \inResetAsync~inputCLKENA0_outclk\ : std_logic;
SIGNAL \GenStrobeI2C|ClkCounter[0]~5_combout\ : std_logic;
SIGNAL \GenStrobeI2C|ClkCounter[0]~DUPLICATE_q\ : std_logic;
SIGNAL \GenStrobeI2C|ClkCounter[1]~4_combout\ : std_logic;
SIGNAL \GenStrobeI2C|ClkCounter[1]~DUPLICATE_q\ : std_logic;
SIGNAL \GenStrobeI2C|ClkCounter[2]~3_combout\ : std_logic;
SIGNAL \GenStrobeI2C|ClkCounter[3]~2_combout\ : std_logic;
SIGNAL \GenStrobeI2C|ClkCounter[4]~1_combout\ : std_logic;
SIGNAL \GenStrobeI2C|ClkCounter[5]~0_combout\ : std_logic;
SIGNAL \GenStrobeI2C|Equal0~0_combout\ : std_logic;
SIGNAL \GenStrobeI2C|oStrobe~q\ : std_logic;
SIGNAL \ConfigureCodec|R.FrameState.Idle~DUPLICATE_q\ : std_logic;
SIGNAL \ConfigureCodec|Add0~25_sumout\ : std_logic;
SIGNAL \ConfigureCodec|Add0~26\ : std_logic;
SIGNAL \ConfigureCodec|Add0~5_sumout\ : std_logic;
SIGNAL \ConfigureCodec|Add0~6\ : std_logic;
SIGNAL \ConfigureCodec|Add0~2\ : std_logic;
SIGNAL \ConfigureCodec|Add0~21_sumout\ : std_logic;
SIGNAL \ConfigureCodec|Add0~22\ : std_logic;
SIGNAL \ConfigureCodec|Add0~17_sumout\ : std_logic;
SIGNAL \ConfigureCodec|Add0~18\ : std_logic;
SIGNAL \ConfigureCodec|Add0~13_sumout\ : std_logic;
SIGNAL \ConfigureCodec|Add0~14\ : std_logic;
SIGNAL \ConfigureCodec|Add0~9_sumout\ : std_logic;
SIGNAL \ConfigureCodec|Equal0~1_combout\ : std_logic;
SIGNAL \ConfigureCodec|Selector1~1_combout\ : std_logic;
SIGNAL \ConfigureCodec|R.FrameState.Start~q\ : std_logic;
SIGNAL \ConfigureCodec|Selector1~0_combout\ : std_logic;
SIGNAL \ConfigureCodec|NextStateAndOutput:vSclkFalling~0_combout\ : std_logic;
SIGNAL \ConfigureCodec|R.BitCtr[3]~DUPLICATE_q\ : std_logic;
SIGNAL \ConfigureCodec|Selector2~0_combout\ : std_logic;
SIGNAL \ConfigureCodec|R.FrameState.Address~q\ : std_logic;
SIGNAL \ConfigureCodec|Selector3~0_combout\ : std_logic;
SIGNAL \ConfigureCodec|R.FrameState.RWBit~q\ : std_logic;
SIGNAL \ConfigureCodec|R.FrameState.Ack1~q\ : std_logic;
SIGNAL \ConfigureCodec|R.FrameState.Ack1~0_combout\ : std_logic;
SIGNAL \ConfigureCodec|R.FrameState.Ack1~DUPLICATE_q\ : std_logic;
SIGNAL \ConfigureCodec|Selector8~0_combout\ : std_logic;
SIGNAL \ConfigureCodec|R.FrameState.Ack3~q\ : std_logic;
SIGNAL \ConfigureCodec|Selector13~0_combout\ : std_logic;
SIGNAL \ioI2cSdin~input_o\ : std_logic;
SIGNAL \ConfigureCodec|Selector16~1_combout\ : std_logic;
SIGNAL \ConfigureCodec|R.AckError~q\ : std_logic;
SIGNAL \ConfigureCodec|Selector5~0_combout\ : std_logic;
SIGNAL \ConfigureCodec|R.FrameState.Data1~q\ : std_logic;
SIGNAL \ConfigureCodec|Selector5~1_combout\ : std_logic;
SIGNAL \ConfigureCodec|R.FrameState.Data1~DUPLICATE_q\ : std_logic;
SIGNAL \ConfigureCodec|Selector13~2_combout\ : std_logic;
SIGNAL \ConfigureCodec|Selector13~1_combout\ : std_logic;
SIGNAL \ConfigureCodec|NextR~10_combout\ : std_logic;
SIGNAL \ConfigureCodec|Selector13~3_combout\ : std_logic;
SIGNAL \ConfigureCodec|Mux8~0_combout\ : std_logic;
SIGNAL \ConfigureCodec|Selector11~2_combout\ : std_logic;
SIGNAL \ConfigureCodec|R.BitCtr[0]~DUPLICATE_q\ : std_logic;
SIGNAL \ConfigureCodec|Selector11~1_combout\ : std_logic;
SIGNAL \ConfigureCodec|Selector11~0_combout\ : std_logic;
SIGNAL \ConfigureCodec|Selector11~3_combout\ : std_logic;
SIGNAL \ConfigureCodec|NextR~8_combout\ : std_logic;
SIGNAL \ConfigureCodec|R.FrameState.Data2~q\ : std_logic;
SIGNAL \ConfigureCodec|Selector7~0_combout\ : std_logic;
SIGNAL \ConfigureCodec|R.FrameState.Data2~DUPLICATE_q\ : std_logic;
SIGNAL \ConfigureCodec|Selector10~0_combout\ : std_logic;
SIGNAL \ConfigureCodec|Selector12~1_combout\ : std_logic;
SIGNAL \ConfigureCodec|Selector12~0_combout\ : std_logic;
SIGNAL \ConfigureCodec|Selector12~2_combout\ : std_logic;
SIGNAL \ConfigureCodec|NextR~9_combout\ : std_logic;
SIGNAL \ConfigureCodec|Selector10~1_combout\ : std_logic;
SIGNAL \ConfigureCodec|Selector10~2_combout\ : std_logic;
SIGNAL \ConfigureCodec|Selector6~0_combout\ : std_logic;
SIGNAL \ConfigureCodec|R.FrameState.Ack2~q\ : std_logic;
SIGNAL \ConfigureCodec|Selector9~0_combout\ : std_logic;
SIGNAL \ConfigureCodec|R.FrameState.Stop~q\ : std_logic;
SIGNAL \ConfigureCodec|R.AddrCtr[6]~1_combout\ : std_logic;
SIGNAL \ConfigureCodec|R.Configured~0_combout\ : std_logic;
SIGNAL \ConfigureCodec|R.Configured~q\ : std_logic;
SIGNAL \WaitCtr[1]~0_combout\ : std_logic;
SIGNAL \WaitCtr[0]~1_combout\ : std_logic;
SIGNAL \WaitCtr[0]~DUPLICATE_q\ : std_logic;
SIGNAL \Start~0_combout\ : std_logic;
SIGNAL \Start~q\ : std_logic;
SIGNAL \ConfigureCodec|R.AddrCtr[6]~0_combout\ : std_logic;
SIGNAL \ConfigureCodec|R.AddrCtr[6]~2_combout\ : std_logic;
SIGNAL \ConfigureCodec|Add0~1_sumout\ : std_logic;
SIGNAL \ConfigureCodec|R.AddrCtr[2]~DUPLICATE_q\ : std_logic;
SIGNAL \ConfigureCodec|R.AddrCtr[1]~DUPLICATE_q\ : std_logic;
SIGNAL \ConfigureCodec|Equal0~0_combout\ : std_logic;
SIGNAL \ConfigureCodec|R.Activity~0_combout\ : std_logic;
SIGNAL \ConfigureCodec|Selector16~0_combout\ : std_logic;
SIGNAL \ConfigureCodec|R.Activity~1_combout\ : std_logic;
SIGNAL \ConfigureCodec|R.Activity~q\ : std_logic;
SIGNAL \ConfigureCodec|Selector0~0_combout\ : std_logic;
SIGNAL \ConfigureCodec|R.FrameState.Idle~q\ : std_logic;
SIGNAL \ConfigureCodec|Selector14~0_combout\ : std_logic;
SIGNAL \ConfigureCodec|R.Sclk~q\ : std_logic;
SIGNAL \ConfigureCodec|Selector15~1_combout\ : std_logic;
SIGNAL \ConfigureCodec|Selector15~2_combout\ : std_logic;
SIGNAL \ConfigureCodec|R.Data[15]~0_combout\ : std_logic;
SIGNAL \ConfigureCodec|Mux0~0_combout\ : std_logic;
SIGNAL \ConfigureCodec|Mux4~0_combout\ : std_logic;
SIGNAL \ConfigureCodec|Mux9~3_combout\ : std_logic;
SIGNAL \ConfigureCodec|Mux6~0_combout\ : std_logic;
SIGNAL \ConfigureCodec|Mux2~0_combout\ : std_logic;
SIGNAL \ConfigureCodec|Mux9~2_combout\ : std_logic;
SIGNAL \ConfigureCodec|Mux5~0_combout\ : std_logic;
SIGNAL \ConfigureCodec|Mux1~0_combout\ : std_logic;
SIGNAL \ConfigureCodec|Mux9~1_combout\ : std_logic;
SIGNAL \ConfigureCodec|Mux3~0_combout\ : std_logic;
SIGNAL \ConfigureCodec|Mux7~0_combout\ : std_logic;
SIGNAL \ConfigureCodec|Mux9~0_combout\ : std_logic;
SIGNAL \ConfigureCodec|Mux9~4_combout\ : std_logic;
SIGNAL \ConfigureCodec|Selector15~0_combout\ : std_logic;
SIGNAL \ConfigureCodec|Selector15~3_combout\ : std_logic;
SIGNAL \ConfigureCodec|R.Sdin~q\ : std_logic;
SIGNAL \iClk~inputCLKENA0_outclk\ : std_logic;
SIGNAL \iSwitch[0]~input_o\ : std_logic;
SIGNAL \ConfigureCodec|R.Configured~DUPLICATE_q\ : std_logic;
SIGNAL \GenClks|Add0~9_sumout\ : std_logic;
SIGNAL \GenClks|ClkCounter[0]~0_combout\ : std_logic;
SIGNAL \GenClks|BMclk~0_combout\ : std_logic;
SIGNAL \GenClks|BMclk~q\ : std_logic;
SIGNAL \GenClks|ADClrc~0_combout\ : std_logic;
SIGNAL \GenClks|Add0~10\ : std_logic;
SIGNAL \GenClks|Add0~5_sumout\ : std_logic;
SIGNAL \GenClks|Add0~6\ : std_logic;
SIGNAL \GenClks|Add0~1_sumout\ : std_logic;
SIGNAL \GenClks|Add0~2\ : std_logic;
SIGNAL \GenClks|Add0~29_sumout\ : std_logic;
SIGNAL \GenClks|BitCounter[1]~DUPLICATE_q\ : std_logic;
SIGNAL \GenClks|BitCounter~1_combout\ : std_logic;
SIGNAL \GenClks|Add0~30\ : std_logic;
SIGNAL \GenClks|Add0~25_sumout\ : std_logic;
SIGNAL \GenClks|Add0~26\ : std_logic;
SIGNAL \GenClks|Add0~21_sumout\ : std_logic;
SIGNAL \GenClks|Add0~22\ : std_logic;
SIGNAL \GenClks|Add0~17_sumout\ : std_logic;
SIGNAL \GenClks|Add0~18\ : std_logic;
SIGNAL \GenClks|Add0~13_sumout\ : std_logic;
SIGNAL \GenClks|BitCounter~0_combout\ : std_logic;
SIGNAL \GenClks|Equal0~0_combout\ : std_logic;
SIGNAL \GenClks|ADClrc~1_combout\ : std_logic;
SIGNAL \GenClks|ADClrc~q\ : std_logic;
SIGNAL \TheI2sToPar|LrcDlyd~q\ : std_logic;
SIGNAL \TheI2sToPar|BclkDlyd~q\ : std_logic;
SIGNAL \TheI2sToPar|BclkRiseEdge~combout\ : std_logic;
SIGNAL \TheI2sToPar|State~0_combout\ : std_logic;
SIGNAL \TheI2sToPar|State~q\ : std_logic;
SIGNAL \TheI2sToPar|NextAudioBitCtr[0]~4_combout\ : std_logic;
SIGNAL \TheI2sToPar|NextAudioBitCtr[1]~3_combout\ : std_logic;
SIGNAL \TheI2sToPar|AudioBitCtr[1]~DUPLICATE_q\ : std_logic;
SIGNAL \TheI2sToPar|NextAudioBitCtr[2]~2_combout\ : std_logic;
SIGNAL \TheI2sToPar|AudioBitCtr[2]~DUPLICATE_q\ : std_logic;
SIGNAL \TheI2sToPar|Equal0~0_combout\ : std_logic;
SIGNAL \TheI2sToPar|NextAudioBitCtr[3]~0_combout\ : std_logic;
SIGNAL \TheI2sToPar|NextAudioBitCtr[4]~1_combout\ : std_logic;
SIGNAL \TheI2sToPar|Equal0~1_combout\ : std_logic;
SIGNAL \TheI2sToPar|NextValL~0_combout\ : std_logic;
SIGNAL \TheI2sToPar|ValL~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[0]~8_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:0:Bandpass0|Add2~34\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:0:Bandpass0|Add2~29_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[1]~7_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[1]~DUPLICATE_q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[0]~DUPLICATE_q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[2]~DUPLICATE_q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:0:Bandpass0|Add2~30\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:0:Bandpass0|Add2~25_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[2]~6_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:11:Bandpass1|Equal1~1_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:0:Bandpass0|Add2~26\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:0:Bandpass0|Add2~21_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[3]~5_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:0:Bandpass0|Add2~22\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:0:Bandpass0|Add2~17_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[4]~4_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:0:Bandpass0|Add2~18\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:0:Bandpass0|Add2~13_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[5]~3_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:0:Bandpass0|Add2~14\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:0:Bandpass0|Add2~9_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[6]~2_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[6]~DUPLICATE_q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[4]~DUPLICATE_q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:0:Bandpass0|Add2~10\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:0:Bandpass0|Add2~5_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[7]~1_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[7]~DUPLICATE_q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:0:Bandpass0|Add2~6\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:0:Bandpass0|Add2~1_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[8]~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[5]~DUPLICATE_q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:11:Bandpass1|Equal1~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:11:Bandpass0|R.SumState.SumValid~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:11:Bandpass0|Selector0~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:11:Bandpass0|R.SumState.Idle~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:11:Bandpass0|Selector1~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:11:Bandpass0|R.SumState.SumEnable~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:11:Bandpass0|Selector2~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:11:Bandpass0|R.SumState.SumSelect~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:11:Bandpass0|Selector3~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:11:Bandpass0|R.SumState.SumWait1~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:11:Bandpass0|R.SumState.SumWait2~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:11:Bandpass0|Selector8~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:11:Bandpass0|R.ValWet~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|R.AddressState~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|R.AddressState~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add2~18\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add2~13_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|R.ReadAddressCoef[1]~3_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add2~14\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add2~25_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|R.ReadAddressCoef[2]~6_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add2~26\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add2~21_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|R.ReadAddressCoef[3]~5_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add2~22\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add2~9_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|R.ReadAddressCoef[4]~2_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add2~10\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add2~5_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|R.ReadAddressCoef[5]~1_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|CoefMemory~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|R.ReadAddressCoef[0]~4_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Equal1~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add2~6\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add2~1_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|R.ReadAddressCoef[6]~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|R.ReadAddressCoef[6]~DUPLICATE_q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|CoefMemory~34_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|CoefMemory~33_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|CoefMemory~35_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|CoefMemory~31_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|CoefMemory~30_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|CoefMemory~32_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|CoefMemory~28_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|CoefMemory~27_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|CoefMemory~29_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|CoefMemory~25_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|CoefMemory~24_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|CoefMemory~26_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|CoefMemory~21_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|CoefMemory~22_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|CoefMemory~23_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|CoefMemory~18_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|CoefMemory~19_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|CoefMemory~20_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|CoefMemory~16_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|CoefMemory~15_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|CoefMemory~17_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|CoefMemory~13_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|CoefMemory~12_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|CoefMemory~14_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|CoefMemory~9_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|CoefMemory~10_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|CoefMemory~11_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|CoefMemory~2_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|CoefMemory~1_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|CoefMemory~3_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|CoefMemory~4_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|CoefMemory~5_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|CoefMemory~6_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|CoefMemory~7_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|CoefMemory~8_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a0~portadataout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a1\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a2\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a3\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a4\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a5\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a6\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a7\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a8\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a9\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a10\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a11\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a12~portadataout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a13\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a14\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a15\ : std_logic;
SIGNAL \iADCdat~input_o\ : std_logic;
SIGNAL \TheI2sToPar|Decoder0~0_combout\ : std_logic;
SIGNAL \TheI2sToPar|D[0]~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-15]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[0]~1_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[0]~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[0]~_wirecell_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add1~2\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add1~5_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add1~6\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add1~9_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add1~10\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add1~13_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add1~14\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add1~17_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add1~18\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add1~21_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add1~22\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add1~25_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add1~26\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add1~29_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add1~30\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add1~33_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[8]~2_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Equal2~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Equal2~1_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[5]~DUPLICATE_q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[8]~_wirecell_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add0~1_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add0~2\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add0~6\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add0~9_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add0~10\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add0~13_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add0~14\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add0~17_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add0~18\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add0~21_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add0~22\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add0~25_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add0~26\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add0~29_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add0~30\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add0~33_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|NextR~7_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Equal0~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add0~5_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|NextR~6_combout\ : std_logic;
SIGNAL \TheI2sToPar|Decoder0~4_combout\ : std_logic;
SIGNAL \TheI2sToPar|D[1]~8_combout\ : std_logic;
SIGNAL \TheI2sToPar|D[2]~2_combout\ : std_logic;
SIGNAL \TheI2sToPar|D[3]~10_combout\ : std_logic;
SIGNAL \TheI2sToPar|Equal0~2_combout\ : std_logic;
SIGNAL \TheI2sToPar|D[4]~4_combout\ : std_logic;
SIGNAL \TheI2sToPar|D[5]~12_combout\ : std_logic;
SIGNAL \TheI2sToPar|Decoder0~3_combout\ : std_logic;
SIGNAL \TheI2sToPar|D[6]~6_combout\ : std_logic;
SIGNAL \TheI2sToPar|D[7]~14_combout\ : std_logic;
SIGNAL \TheI2sToPar|Decoder0~1_combout\ : std_logic;
SIGNAL \TheI2sToPar|D[8]~1_combout\ : std_logic;
SIGNAL \TheI2sToPar|D[9]~9_combout\ : std_logic;
SIGNAL \TheI2sToPar|D[10]~3_combout\ : std_logic;
SIGNAL \TheI2sToPar|D[11]~11_combout\ : std_logic;
SIGNAL \TheI2sToPar|Decoder0~2_combout\ : std_logic;
SIGNAL \TheI2sToPar|D[12]~5_combout\ : std_logic;
SIGNAL \TheI2sToPar|D[13]~13_combout\ : std_logic;
SIGNAL \TheI2sToPar|D[14]~7_combout\ : std_logic;
SIGNAL \TheI2sToPar|D[14]~feeder_combout\ : std_logic;
SIGNAL \TheI2sToPar|D[15]~15_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a0~portbdataout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-15]~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-14]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a1\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-14]~1_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-13]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a2\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-13]~2_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-12]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a3\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-12]~3_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-11]~feeder_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-11]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a4\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-11]~4_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a5\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-10]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-10]~5_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-9]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a6\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-9]~6_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-8]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a7\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-8]~7_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-7]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a8\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-7]~8_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-6]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a9\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-6]~9_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a10\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-5]~feeder_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-5]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-5]~10_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-4]~feeder_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-4]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a11\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-4]~11_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-3]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a12~portbdataout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-3]~12_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-2]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a13\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-2]~13_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a14\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-1]~feeder_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-1]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-1]~14_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[0]~DUPLICATE_q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a15\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Sample[0]~15_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~39\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~38\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~37\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~36\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~35\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~34\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~33\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~32\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~31\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~30\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~29\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~28\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~27\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~26\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~25\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~24\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~19\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~20\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~22\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~12\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~10\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~11\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~21\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_resulta\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|vAdd~2_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~13\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~14\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~16\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~15\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~18\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~17\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~9\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|vAdd~1_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|vAdd~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~23\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add3~14\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add3~18\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add3~22\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add3~26\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add3~30\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add3~34\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add3~38\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add3~42\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add3~46\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add3~50\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add3~54\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add3~58\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add3~62\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add3~66\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add3~70\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add3~10\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add3~6\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add3~1_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[0]~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add3~9_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM77\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add3~69_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-1]_OTERM99\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add3~5_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM75\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM73\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-1]~14_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add3~65_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-2]_OTERM105\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-2]~13_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add3~61_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-3]_OTERM111\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-3]~12_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add3~57_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-4]_OTERM117\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-4]~11_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add3~53_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-5]_OTERM123\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-5]~10_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add3~49_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-6]_OTERM129\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-6]~9_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add3~45_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-7]_OTERM135\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-7]~8_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add3~41_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-8]_OTERM141\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-8]~7_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add3~37_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-9]_OTERM147\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-9]~6_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add3~33_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-10]_OTERM153\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-10]~5_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add3~29_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-11]_OTERM159\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-11]~4_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add3~25_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-12]_OTERM165\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-12]~3_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add3~21_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-13]_OTERM171\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-13]~2_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add3~17_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-14]_OTERM177\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-14]~1_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add3~13_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM79\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-15]~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add4~5_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-15]~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Selector2~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|R.SumState.SumSelect~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Selector3~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|R.SumState.SumWait1~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|R.SumState.SumWait2~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|R.SumState.SumValid~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Selector0~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|R.SumState.Idle~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Selector1~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|R.SumState.SumEnable~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Selector6~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|R.SelSumUp~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Selector7~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|R.EnableSumUp~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-15]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add4~10\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add4~13_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-14]~1_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-14]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add4~14\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add4~17_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-13]~2_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-13]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add4~18\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add4~21_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-12]~3_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-12]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add4~22\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add4~25_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-11]~4_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-11]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add4~26\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add4~29_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-10]~5_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-10]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add4~30\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add4~33_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-9]~6_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-9]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add4~34\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add4~37_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-8]~7_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-8]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add4~38\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add4~41_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-7]~8_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-7]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add4~42\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add4~45_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-6]~9_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-6]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add4~46\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add4~49_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-5]~10_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-5]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add4~50\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add4~53_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-4]~11_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-4]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add4~54\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add4~57_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-3]~12_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-3]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add4~58\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add4~61_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-2]~13_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-2]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add4~62\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add4~65_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-1]~14_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-1]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add4~66\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add4~6\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add4~1_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Add4~1_wirecell_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a0\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a1\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a2\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a3\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a4\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a5\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a6\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a7\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a8\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a9\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a10\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a11\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a12\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a13\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a14\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a15\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a0\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-15]~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a1\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-14]~1_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a2\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-13]~2_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a3\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-12]~3_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a4\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-11]~4_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a5\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-10]~5_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a6\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-9]~6_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a7\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-8]~7_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a8\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-7]~8_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a9\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-6]~9_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a10\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-5]~10_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a11\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-4]~11_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a12\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-3]~12_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a13\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-2]~13_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a14\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-1]~14_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a15\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Sample[0]~15_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~39\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~38\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~37\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~36\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~35\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~34\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~33\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~32\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~31\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~30\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~29\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~28\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~27\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~26\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~25\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~24\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~23\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~16\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~18\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~17\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~15\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~14\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~9\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|vAdd~1_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~20\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~22\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~13\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~12\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_resulta\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~21\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~10\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~11\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|vAdd~2_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~19\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|vAdd~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add3~14\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add3~18\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add3~22\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add3~26\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add3~30\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add3~34\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add3~38\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add3~42\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add3~46\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add3~50\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add3~54\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add3~58\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add3~62\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add3~66\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add3~70\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add3~10\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add3~6\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add3~1_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[0]~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add3~9_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM69\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add3~69_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-1]_OTERM97\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add3~5_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM67\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM65\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-1]~14_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add3~65_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-2]_OTERM103\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-2]~13_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add4~5_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add3~61_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-3]_OTERM109\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-3]~12_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add3~57_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-4]_OTERM115\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-4]~11_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add3~53_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-5]_OTERM121\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-5]~10_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add3~49_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-6]_OTERM127\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-6]~9_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add3~45_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-7]_OTERM133\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-7]~8_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add3~41_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-8]_OTERM139\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-8]~7_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add3~37_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-9]_OTERM145\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-9]~6_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add3~33_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-10]_OTERM151\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-10]~5_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add3~29_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-11]_OTERM157\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-11]~4_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add3~25_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-12]_OTERM163\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-12]~3_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add3~21_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-13]_OTERM169\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-13]~2_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add3~17_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-14]_OTERM175\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-14]~1_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add3~13_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM71\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-15]~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-15]~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|R.SumState.SumValid~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Selector0~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|R.SumState.Idle~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Selector1~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|R.SumState.SumEnable~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Selector2~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|R.SumState.SumSelect~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Selector3~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|R.SumState.SumWait1~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|R.SumState.SumWait2~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Selector6~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|R.SelSumUp~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|R.SumState.Idle~DUPLICATE_q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Selector7~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|R.EnableSumUp~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-15]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add4~10\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add4~13_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-14]~1_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-14]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add4~14\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add4~17_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-13]~2_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-13]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add4~18\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add4~21_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-12]~3_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-12]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add4~22\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add4~25_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-11]~4_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-11]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add4~26\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add4~29_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-10]~5_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-10]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add4~30\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add4~33_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-9]~6_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-9]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add4~34\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add4~37_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-8]~7_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-8]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add4~38\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add4~41_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-7]~8_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-7]~DUPLICATE_q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add4~42\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add4~45_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-6]~9_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-6]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add4~46\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add4~49_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-5]~10_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-5]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add4~50\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add4~53_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-4]~11_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-4]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add4~54\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add4~57_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-3]~12_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-3]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add4~58\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add4~61_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-2]~13_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-2]~DUPLICATE_q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add4~62\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add4~65_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-1]~14_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-1]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add4~66\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add4~6\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add4~1_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Add4~1_wirecell_combout\ : std_logic;
SIGNAL \TheRxFsk|Mux1~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-2]~q\ : std_logic;
SIGNAL \TheRxFsk|Mux2~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-3]~DUPLICATE_q\ : std_logic;
SIGNAL \TheRxFsk|Mux3~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-4]~DUPLICATE_q\ : std_logic;
SIGNAL \TheRxFsk|Mux4~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Mux5~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Mux6~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-7]~q\ : std_logic;
SIGNAL \TheRxFsk|Mux7~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-8]~DUPLICATE_q\ : std_logic;
SIGNAL \TheRxFsk|Mux8~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Mux9~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Mux10~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Mux11~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Mux12~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Mux13~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Mux14~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Mux15~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Add0~6\ : std_logic;
SIGNAL \TheRxFsk|Add0~10\ : std_logic;
SIGNAL \TheRxFsk|Add0~14\ : std_logic;
SIGNAL \TheRxFsk|Add0~18\ : std_logic;
SIGNAL \TheRxFsk|Add0~22\ : std_logic;
SIGNAL \TheRxFsk|Add0~26\ : std_logic;
SIGNAL \TheRxFsk|Add0~30\ : std_logic;
SIGNAL \TheRxFsk|Add0~34\ : std_logic;
SIGNAL \TheRxFsk|Add0~38\ : std_logic;
SIGNAL \TheRxFsk|Add0~42\ : std_logic;
SIGNAL \TheRxFsk|Add0~46\ : std_logic;
SIGNAL \TheRxFsk|Add0~50\ : std_logic;
SIGNAL \TheRxFsk|Add0~54\ : std_logic;
SIGNAL \TheRxFsk|Add0~58\ : std_logic;
SIGNAL \TheRxFsk|Add0~62\ : std_logic;
SIGNAL \TheRxFsk|Add0~1_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a0~portadataout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a1\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a2\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a3\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a4~portadataout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a5\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a6\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a7\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a8\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a9\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a10\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a11\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a12\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a13\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a14\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a15\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a0~portbdataout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-15]~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a1\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-14]~1_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a2\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-13]~2_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a3\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-12]~3_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a4~portbdataout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-11]~4_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a5\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-10]~5_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a6\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-9]~6_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a7\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-8]~7_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a8\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-7]~8_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a9\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-6]~9_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a10\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-5]~10_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a11\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-4]~11_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a12\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-3]~12_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a13\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-2]~13_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a14\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-1]~14_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a15\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Sample[0]~15_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~39\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~38\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~37\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~36\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~35\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~34\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~33\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~32\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~31\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~30\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~29\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~28\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~27\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~26\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~25\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~24\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~23\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~20\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~22\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~13\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~19\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~21\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~10\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~11\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~12\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_resulta\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|vAdd~2_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~15\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~18\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~17\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~16\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~14\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~9\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|vAdd~1_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|vAdd~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add3~14\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add3~18\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add3~22\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add3~26\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add3~30\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add3~34\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add3~38\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add3~42\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add3~46\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add3~50\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add3~54\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add3~58\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add3~62\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add3~66\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add3~70\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add3~10\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add3~6\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add3~1_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[0]~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add3~9_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM85\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM81\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add3~5_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM83\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add3~69_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-1]_OTERM101\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-1]~14_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add3~65_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-2]_OTERM107\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-2]~13_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add4~5_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add3~61_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-3]_OTERM113\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-3]~12_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add3~57_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-4]_OTERM119\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-4]~11_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add3~53_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-5]_OTERM125\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-5]~10_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add3~49_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-6]_OTERM131\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-6]~9_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add3~45_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-7]_OTERM137\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-7]~8_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add3~41_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-8]_OTERM143\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-8]~7_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add3~37_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-9]_OTERM149\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-9]~6_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add3~33_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-10]_OTERM155\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-10]~5_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add3~29_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-11]_OTERM161\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-11]~4_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add3~25_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-12]_OTERM167\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-12]~3_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add3~21_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-13]_OTERM173\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-13]~2_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add3~17_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-14]_OTERM179\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-14]~1_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add3~13_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM87\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-15]~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-15]~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|R.SumState.SumValid~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Selector0~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|R.SumState.Idle~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Selector1~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|R.SumState.SumEnable~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Selector2~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|R.SumState.SumSelect~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Selector3~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|R.SumState.SumWait1~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|R.SumState.SumWait2~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Selector6~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|R.SelSumUp~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Selector7~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|R.EnableSumUp~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-15]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add4~10\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add4~13_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-14]~1_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-14]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add4~14\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add4~17_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-13]~2_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-13]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add4~18\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add4~21_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-12]~3_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-12]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add4~22\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add4~25_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-11]~4_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-11]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add4~26\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add4~29_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-10]~5_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-10]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add4~30\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add4~33_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-9]~6_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-9]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add4~34\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add4~37_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-8]~7_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-8]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add4~38\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add4~41_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-7]~8_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-7]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add4~42\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add4~45_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-6]~9_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-6]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add4~46\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add4~49_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-5]~10_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-5]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add4~50\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add4~53_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-4]~11_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-4]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add4~54\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add4~57_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-3]~12_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-3]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add4~58\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add4~61_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-2]~13_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-2]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add4~62\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add4~65_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-1]~14_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-1]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add4~66\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add4~6\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add4~1_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Add4~1_wirecell_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a0\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a1\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a2\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a3\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a4\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a5\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a6\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a7\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a8\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a9\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a10\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a11\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a12\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a13\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a14\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a15\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a0\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-15]~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a1\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-14]~1_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a2\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-13]~2_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a3\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-12]~3_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a4\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-11]~4_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a5\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-10]~5_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a6\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-9]~6_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a7\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-8]~7_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a8\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-7]~8_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a9\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-6]~9_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a10\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-5]~10_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a11\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-4]~11_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a12\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-3]~12_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a13\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-2]~13_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a14\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-1]~14_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a15\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Sample[0]~15_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~39\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~38\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~37\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~36\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~35\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~34\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~33\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~32\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~31\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~30\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~29\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~28\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~27\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~26\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~25\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~24\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~23\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~19\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~15\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~18\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~17\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~16\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~14\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~9\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|vAdd~1_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~22\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~20\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~13\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~11\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~12\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~21\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~10\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_resulta\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|vAdd~2_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|vAdd~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add3~14\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add3~18\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add3~22\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add3~26\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add3~30\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add3~34\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add3~38\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add3~42\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add3~46\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add3~50\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add3~54\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add3~58\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add3~62\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add3~66\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add3~70\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add3~10\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add3~6\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add3~1_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[0]~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add3~9_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM13\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add3~5_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM11\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM9\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add3~69_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-1]_OTERM17\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-1]~14_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add4~5_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add3~65_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-2]_OTERM21\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-2]~13_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add3~61_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-3]_OTERM25\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-3]~12_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add3~57_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-4]_OTERM29\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-4]~11_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add3~53_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-5]_OTERM33\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-5]~10_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add3~49_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-6]_OTERM37\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-6]~9_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add3~45_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-7]_OTERM43\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-7]~8_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add3~41_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-8]_OTERM47\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-8]~7_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add3~37_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-9]_OTERM53\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-9]~6_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add3~33_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-10]_OTERM55\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-10]~5_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add3~29_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-11]_OTERM59\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-11]~4_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add3~25_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-12]_OTERM63\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-12]~3_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add3~21_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-13]_OTERM91\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-13]~2_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add3~17_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-14]_OTERM95\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-14]~1_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add3~13_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM15\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-15]~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-15]~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|R.SumState.SumEnable~DUPLICATE_q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Selector2~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|R.SumState.SumSelect~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Selector3~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|R.SumState.SumWait1~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|R.SumState.SumWait2~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|R.SumState.SumValid~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Selector0~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|R.SumState.Idle~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Selector1~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|R.SumState.SumEnable~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Selector6~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|R.SelSumUp~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Selector7~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|R.EnableSumUp~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-15]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add4~10\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add4~13_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-14]~1_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-14]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add4~14\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add4~17_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-13]~2_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-13]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add4~18\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add4~21_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-12]~3_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-12]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add4~22\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add4~25_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-11]~4_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-11]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add4~26\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add4~29_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-10]~5_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-10]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add4~30\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add4~33_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-9]~6_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-9]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add4~34\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add4~37_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-8]~7_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-8]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add4~38\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add4~41_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-7]~8_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-7]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add4~42\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add4~45_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-6]~9_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-6]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add4~46\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add4~49_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-5]~10_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-5]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add4~50\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add4~53_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-4]~11_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-4]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add4~54\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add4~57_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-3]~12_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-3]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add4~58\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add4~61_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-2]~13_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-2]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add4~62\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add4~65_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-1]~14_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-1]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add4~66\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add4~6\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add4~1_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Add4~1_wirecell_combout\ : std_logic;
SIGNAL \TheRxFsk|Mux17~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Mux18~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-3]~DUPLICATE_q\ : std_logic;
SIGNAL \TheRxFsk|Mux19~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Mux20~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Mux21~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Mux22~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Mux23~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Mux24~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Mux25~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Mux26~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Mux27~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Mux28~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Mux29~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Mux30~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Mux31~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Add1~6\ : std_logic;
SIGNAL \TheRxFsk|Add1~10\ : std_logic;
SIGNAL \TheRxFsk|Add1~14\ : std_logic;
SIGNAL \TheRxFsk|Add1~18\ : std_logic;
SIGNAL \TheRxFsk|Add1~22\ : std_logic;
SIGNAL \TheRxFsk|Add1~26\ : std_logic;
SIGNAL \TheRxFsk|Add1~30\ : std_logic;
SIGNAL \TheRxFsk|Add1~34\ : std_logic;
SIGNAL \TheRxFsk|Add1~38\ : std_logic;
SIGNAL \TheRxFsk|Add1~42\ : std_logic;
SIGNAL \TheRxFsk|Add1~46\ : std_logic;
SIGNAL \TheRxFsk|Add1~50\ : std_logic;
SIGNAL \TheRxFsk|Add1~54\ : std_logic;
SIGNAL \TheRxFsk|Add1~58\ : std_logic;
SIGNAL \TheRxFsk|Add1~62\ : std_logic;
SIGNAL \TheRxFsk|Add1~1_sumout\ : std_logic;
SIGNAL \TheRxFsk|Add0~61_sumout\ : std_logic;
SIGNAL \TheRxFsk|Add1~61_sumout\ : std_logic;
SIGNAL \TheRxFsk|Add1~57_sumout\ : std_logic;
SIGNAL \TheRxFsk|Add0~57_sumout\ : std_logic;
SIGNAL \TheRxFsk|Add0~53_sumout\ : std_logic;
SIGNAL \TheRxFsk|Add1~53_sumout\ : std_logic;
SIGNAL \TheRxFsk|Add1~49_sumout\ : std_logic;
SIGNAL \TheRxFsk|Add0~49_sumout\ : std_logic;
SIGNAL \TheRxFsk|Add1~45_sumout\ : std_logic;
SIGNAL \TheRxFsk|Add0~45_sumout\ : std_logic;
SIGNAL \TheRxFsk|Add0~41_sumout\ : std_logic;
SIGNAL \TheRxFsk|Add1~41_sumout\ : std_logic;
SIGNAL \TheRxFsk|Add1~37_sumout\ : std_logic;
SIGNAL \TheRxFsk|Add0~37_sumout\ : std_logic;
SIGNAL \TheRxFsk|Add1~33_sumout\ : std_logic;
SIGNAL \TheRxFsk|Add0~33_sumout\ : std_logic;
SIGNAL \TheRxFsk|Add1~29_sumout\ : std_logic;
SIGNAL \TheRxFsk|Add0~29_sumout\ : std_logic;
SIGNAL \TheRxFsk|Add1~25_sumout\ : std_logic;
SIGNAL \TheRxFsk|Add0~25_sumout\ : std_logic;
SIGNAL \TheRxFsk|Add1~21_sumout\ : std_logic;
SIGNAL \TheRxFsk|Add0~21_sumout\ : std_logic;
SIGNAL \TheRxFsk|Add1~17_sumout\ : std_logic;
SIGNAL \TheRxFsk|Add0~17_sumout\ : std_logic;
SIGNAL \TheRxFsk|Add1~13_sumout\ : std_logic;
SIGNAL \TheRxFsk|Add0~13_sumout\ : std_logic;
SIGNAL \TheRxFsk|Add1~9_sumout\ : std_logic;
SIGNAL \TheRxFsk|Add0~9_sumout\ : std_logic;
SIGNAL \TheRxFsk|Add1~5_sumout\ : std_logic;
SIGNAL \TheRxFsk|Add0~5_sumout\ : std_logic;
SIGNAL \TheRxFsk|Add2~70_cout\ : std_logic;
SIGNAL \TheRxFsk|Add2~10\ : std_logic;
SIGNAL \TheRxFsk|Add2~14\ : std_logic;
SIGNAL \TheRxFsk|Add2~18\ : std_logic;
SIGNAL \TheRxFsk|Add2~22\ : std_logic;
SIGNAL \TheRxFsk|Add2~26\ : std_logic;
SIGNAL \TheRxFsk|Add2~30\ : std_logic;
SIGNAL \TheRxFsk|Add2~34\ : std_logic;
SIGNAL \TheRxFsk|Add2~38\ : std_logic;
SIGNAL \TheRxFsk|Add2~42\ : std_logic;
SIGNAL \TheRxFsk|Add2~46\ : std_logic;
SIGNAL \TheRxFsk|Add2~50\ : std_logic;
SIGNAL \TheRxFsk|Add2~54\ : std_logic;
SIGNAL \TheRxFsk|Add2~58\ : std_logic;
SIGNAL \TheRxFsk|Add2~62\ : std_logic;
SIGNAL \TheRxFsk|Add2~66\ : std_logic;
SIGNAL \TheRxFsk|Add2~2\ : std_logic;
SIGNAL \TheRxFsk|Add2~5_sumout\ : std_logic;
SIGNAL \TheRxFsk|Add2~1_sumout\ : std_logic;
SIGNAL \TheRxFsk|Add2~9_sumout\ : std_logic;
SIGNAL \TheRxFsk|Substracted[-15]~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|R.WriteAddress[0]~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add1~2\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add1~5_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|R.WriteAddress[1]~1_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add1~6\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add1~9_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|vNextWriteAddress~1_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add1~10\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add1~13_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|R.WriteAddress[3]~2_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add1~14\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add1~17_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|vNextWriteAddress~2_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add1~18\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add1~21_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|vNextWriteAddress~3_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add1~22\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add1~25_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|R.WriteAddress[6]~3_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Equal2~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|vNextWriteAddress~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|R.WriteAddress[0]~DUPLICATE_q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|R.WriteAddress[1]~DUPLICATE_q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|R.WriteAddress[1]~_wirecell_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|R.WriteAddress[3]~_wirecell_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|R.WriteAddress[6]~_wirecell_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add0~2\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add0~5_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add0~6\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add0~9_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add0~10\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add0~13_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|NextR~8_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add0~14\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add0~17_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add0~18\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add0~21_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add0~22\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add0~25_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|NextR~9_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Equal0~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|NextR~7_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|NextR~6_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|R.ReadAddressSample[0]~DUPLICATE_q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|R.ReadAddressSample[1]~DUPLICATE_q\ : std_logic;
SIGNAL \TheRxFsk|Add2~13_sumout\ : std_logic;
SIGNAL \TheRxFsk|Substracted[-14]~1_combout\ : std_logic;
SIGNAL \TheRxFsk|Add2~17_sumout\ : std_logic;
SIGNAL \TheRxFsk|Substracted[-13]~2_combout\ : std_logic;
SIGNAL \TheRxFsk|Add2~21_sumout\ : std_logic;
SIGNAL \TheRxFsk|Substracted[-12]~3_combout\ : std_logic;
SIGNAL \TheRxFsk|Add2~25_sumout\ : std_logic;
SIGNAL \TheRxFsk|Substracted[-11]~4_combout\ : std_logic;
SIGNAL \TheRxFsk|Add2~29_sumout\ : std_logic;
SIGNAL \TheRxFsk|Substracted[-10]~5_combout\ : std_logic;
SIGNAL \TheRxFsk|Add2~33_sumout\ : std_logic;
SIGNAL \TheRxFsk|Substracted[-9]~6_combout\ : std_logic;
SIGNAL \TheRxFsk|Add2~37_sumout\ : std_logic;
SIGNAL \TheRxFsk|Substracted[-8]~7_combout\ : std_logic;
SIGNAL \TheRxFsk|Add2~41_sumout\ : std_logic;
SIGNAL \TheRxFsk|Substracted[-7]~8_combout\ : std_logic;
SIGNAL \TheRxFsk|Add2~45_sumout\ : std_logic;
SIGNAL \TheRxFsk|Substracted[-6]~9_combout\ : std_logic;
SIGNAL \TheRxFsk|Add2~49_sumout\ : std_logic;
SIGNAL \TheRxFsk|Substracted[-5]~10_combout\ : std_logic;
SIGNAL \TheRxFsk|Add2~53_sumout\ : std_logic;
SIGNAL \TheRxFsk|Substracted[-4]~11_combout\ : std_logic;
SIGNAL \TheRxFsk|Add2~57_sumout\ : std_logic;
SIGNAL \TheRxFsk|Substracted[-3]~12_combout\ : std_logic;
SIGNAL \TheRxFsk|Add2~61_sumout\ : std_logic;
SIGNAL \TheRxFsk|Substracted[-2]~13_combout\ : std_logic;
SIGNAL \TheRxFsk|Add2~65_sumout\ : std_logic;
SIGNAL \TheRxFsk|Substracted[-1]~14_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a0~portbdataout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|R.FirstSample~q\ : std_logic;
SIGNAL \TheRxFsk|Add2~5_wirecell_combout\ : std_logic;
SIGNAL \TheRxFsk|result~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|DdryDelayed[-15]~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Sample[-15]~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|DdryDelayed[-14]~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a1\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Sample[-14]~1_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|DdryDelayed[-13]~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a2\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Sample[-13]~2_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a3\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|DdryDelayed[-12]~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Sample[-12]~3_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|DdryDelayed[-11]~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a4\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Sample[-11]~4_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a5\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|DdryDelayed[-10]~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Sample[-10]~5_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|DdryDelayed[-9]~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a6\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Sample[-9]~6_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|DdryDelayed[-8]~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a7\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Sample[-8]~7_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|DdryDelayed[-7]~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a8\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Sample[-7]~8_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a9\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|DdryDelayed[-6]~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Sample[-6]~9_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|DdryDelayed[-5]~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a10\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Sample[-5]~10_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|DdryDelayed[-4]~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a11\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Sample[-4]~11_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a12\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|DdryDelayed[-3]~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Sample[-3]~12_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|DdryDelayed[-2]~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a13\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Sample[-2]~13_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|DdryDelayed[-1]~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a14\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Sample[-1]~14_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a15\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Sample[0]~15_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~39\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~38\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~37\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~36\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~35\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~34\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~33\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~32\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~31\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~30\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~29\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~28\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~27\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~26\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~25\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~24\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~23\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~19\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~17\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~9\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~15\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~16\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~18\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~14\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|vAdd~1_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~8_resulta\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~21\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~10\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~11\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~12\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|vAdd~2_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~22\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~20\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Mult0~13\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|vAdd~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add3~70\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add3~66\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add3~62\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add3~58\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add3~54\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add3~50\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add3~46\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add3~42\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add3~38\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add3~34\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add3~30\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add3~26\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add3~22\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add3~18\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add3~14\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add3~10\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add3~6\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add3~1_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|MultResultDelayed[0]~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add3~9_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM5\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add3~13_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|MultResultDelayed[-1]_OTERM19\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM1\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add3~5_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM3\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|MultResult[-1]~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add4~5_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add3~17_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|MultResultDelayed[-2]_OTERM23\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|MultResult[-2]~1_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add3~21_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|MultResultDelayed[-3]_OTERM27\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|MultResult[-3]~2_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add3~25_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|MultResultDelayed[-4]_OTERM31\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|MultResult[-4]~3_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add3~29_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|MultResultDelayed[-5]_OTERM35\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|MultResult[-5]~4_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add3~33_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|MultResultDelayed[-6]_OTERM39\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|MultResult[-6]~5_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add3~37_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|MultResultDelayed[-7]_OTERM41\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|MultResult[-7]~6_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add3~41_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|MultResultDelayed[-8]_OTERM45\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|MultResult[-8]~7_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add3~45_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|MultResultDelayed[-9]_OTERM51\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|MultResult[-9]~8_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add3~49_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|MultResultDelayed[-10]_OTERM49\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|MultResult[-10]~9_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add3~53_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|MultResultDelayed[-11]_OTERM57\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|MultResult[-11]~10_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add3~57_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|MultResultDelayed[-12]_OTERM61\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|MultResult[-12]~11_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add3~61_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|MultResultDelayed[-13]_OTERM89\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|MultResult[-13]~12_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add3~65_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|MultResultDelayed[-14]_OTERM93\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|MultResult[-14]~13_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add3~69_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM7\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|MultResult[-15]~14_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|NextSum[-15]~14_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|R.SumState.SumValid~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Selector0~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|R.SumState.Idle~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Selector1~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|R.SumState.SumEnable~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Selector2~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|R.SumState.SumSelect~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Selector3~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|R.SumState.SumWait1~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|R.SumState.SumWait2~DUPLICATE_q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Selector6~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|R.SelSumUp~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|R.SumState.SumWait2~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Selector7~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|R.EnableSumUp~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Sum[-15]~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add4~66\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add4~61_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|NextSum[-14]~13_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Sum[-14]~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add4~62\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add4~57_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|NextSum[-13]~12_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Sum[-13]~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add4~58\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add4~53_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|NextSum[-12]~11_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Sum[-12]~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add4~54\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add4~49_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|NextSum[-11]~10_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Sum[-11]~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add4~50\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add4~45_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|NextSum[-10]~9_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Sum[-10]~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add4~46\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add4~41_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|NextSum[-9]~8_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Sum[-9]~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add4~42\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add4~37_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|NextSum[-8]~7_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Sum[-8]~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add4~38\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add4~33_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|NextSum[-7]~6_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Sum[-7]~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add4~34\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add4~29_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|NextSum[-6]~5_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Sum[-6]~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add4~30\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add4~25_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|NextSum[-5]~4_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Sum[-5]~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add4~26\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add4~21_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|NextSum[-4]~3_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Sum[-4]~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add4~22\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add4~17_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|NextSum[-3]~2_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Sum[-3]~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add4~18\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add4~13_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|NextSum[-2]~1_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Sum[-2]~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add4~14\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add4~9_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|NextSum[-1]~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Sum[-1]~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add4~10\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add4~6\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add4~1_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Add4~1_wirecell_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|Selector8~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|R.ValWet~q\ : std_logic;
SIGNAL \TheRxFsk|oD~0_combout\ : std_logic;
SIGNAL \TheRxFsk|oD~q\ : std_logic;
SIGNAL \TheParToI2s|Selector0~0_combout\ : std_logic;
SIGNAL \TheParToI2s|State.WaitingValL~q\ : std_logic;
SIGNAL \TheParToI2s|Selector1~0_combout\ : std_logic;
SIGNAL \TheParToI2s|State.SyncingToBclk~q\ : std_logic;
SIGNAL \TheParToI2s|State.FirstBitEmptyL~0_combout\ : std_logic;
SIGNAL \TheParToI2s|State.FirstBitEmptyL~q\ : std_logic;
SIGNAL \TheParToI2s|Selector3~0_combout\ : std_logic;
SIGNAL \TheParToI2s|State.SendingL~q\ : std_logic;
SIGNAL \TheParToI2s|Selector4~0_combout\ : std_logic;
SIGNAL \TheParToI2s|State.FirstBitEmptyR~q\ : std_logic;
SIGNAL \TheParToI2s|Selector8~0_combout\ : std_logic;
SIGNAL \TheParToI2s|State.SyncingToBclk~DUPLICATE_q\ : std_logic;
SIGNAL \TheParToI2s|NextBclkCtr~0_combout\ : std_logic;
SIGNAL \TheParToI2s|Selector7~0_combout\ : std_logic;
SIGNAL \TheParToI2s|Selector9~0_combout\ : std_logic;
SIGNAL \TheParToI2s|Selector9~1_combout\ : std_logic;
SIGNAL \TheParToI2s|Add0~0_combout\ : std_logic;
SIGNAL \TheParToI2s|Selector7~1_combout\ : std_logic;
SIGNAL \TheParToI2s|NextBclkCtr~1_combout\ : std_logic;
SIGNAL \TheParToI2s|Selector8~1_combout\ : std_logic;
SIGNAL \TheParToI2s|NextState~6_combout\ : std_logic;
SIGNAL \TheParToI2s|Selector5~0_combout\ : std_logic;
SIGNAL \TheParToI2s|State.SendingR~q\ : std_logic;
SIGNAL \TheParToI2s|Selector10~0_combout\ : std_logic;
SIGNAL \TheParToI2s|Selector6~1_combout\ : std_logic;
SIGNAL \TheParToI2s|Selector6~0_combout\ : std_logic;
SIGNAL \TheParToI2s|Selector6~2_combout\ : std_logic;
SIGNAL \TheParToI2s|BclkCtr[3]~DUPLICATE_q\ : std_logic;
SIGNAL \TheParToI2s|LastValidDL[6]~feeder_combout\ : std_logic;
SIGNAL \TheParToI2s|LastValidDL[12]~feeder_combout\ : std_logic;
SIGNAL \TheParToI2s|Mux1~1_combout\ : std_logic;
SIGNAL \TheParToI2s|BclkCtr[2]~DUPLICATE_q\ : std_logic;
SIGNAL \TheParToI2s|Mux1~2_combout\ : std_logic;
SIGNAL \TheParToI2s|LastValidDL[5]~feeder_combout\ : std_logic;
SIGNAL \TheParToI2s|Mux1~3_combout\ : std_logic;
SIGNAL \TheParToI2s|LastValidDL[0]~feeder_combout\ : std_logic;
SIGNAL \TheParToI2s|LastValidDL[8]~feeder_combout\ : std_logic;
SIGNAL \TheParToI2s|Mux1~0_combout\ : std_logic;
SIGNAL \TheParToI2s|Selector10~1_combout\ : std_logic;
SIGNAL \TheParToI2s|oLrc~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\ : std_logic_vector(8 DOWNTO 0);
SIGNAL \TheI2sToPar|AudioBitCtr\ : std_logic_vector(4 DOWNTO 0);
SIGNAL \ConfigureCodec|R.AddrCtr\ : std_logic_vector(6 DOWNTO 0);
SIGNAL \SyncSwitchInput|Metastable\ : std_logic_vector(1 DOWNTO 0);
SIGNAL \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire\ : std_logic_vector(0 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|Sum\ : std_logic_vector(0 DOWNTO 0);
SIGNAL \TheRxFsk|Lowpass|DdryDelayed\ : std_logic_vector(0 DOWNTO 0);
SIGNAL \TheRxFsk|Lowpass|Sum\ : std_logic_vector(0 DOWNTO 0);
SIGNAL \ConfigureCodec|R.BitCtr\ : std_logic_vector(3 DOWNTO 0);
SIGNAL \TheI2sToPar|D\ : std_logic_vector(16 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|Sum\ : std_logic_vector(0 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|Sum\ : std_logic_vector(0 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|Sum\ : std_logic_vector(0 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\ : std_logic_vector(8 DOWNTO 0);
SIGNAL \GenClks|ClkCounter\ : std_logic_vector(0 DOWNTO 0);
SIGNAL \TheParToI2s|LastValidDL\ : std_logic_vector(15 DOWNTO 0);
SIGNAL \GenClks|BitCounter\ : std_logic_vector(7 DOWNTO 0);
SIGNAL \TheParToI2s|BclkCtr\ : std_logic_vector(3 DOWNTO 0);
SIGNAL WaitCtr : std_logic_vector(1 DOWNTO 0);
SIGNAL \GenStrobeI2C|ClkCounter\ : std_logic_vector(5 DOWNTO 0);
SIGNAL \TheRxFsk|Lowpass|MultResultDelayed\ : std_logic_vector(0 DOWNTO 0);
SIGNAL \ConfigureCodec|R.Data\ : std_logic_vector(15 DOWNTO 0);
SIGNAL \TheRxFsk|Lowpass|R.ReadAddressCoef\ : std_logic_vector(6 DOWNTO 0);
SIGNAL \TheRxFsk|Lowpass|R.WriteAddress\ : std_logic_vector(6 DOWNTO 0);
SIGNAL \TheRxFsk|Lowpass|R.ReadAddressSample\ : std_logic_vector(6 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed\ : std_logic_vector(0 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed\ : std_logic_vector(0 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed\ : std_logic_vector(0 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed\ : std_logic_vector(0 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed\ : std_logic_vector(0 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\ : std_logic_vector(8 DOWNTO 0);
SIGNAL \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|fboutclk_wire\ : std_logic_vector(0 DOWNTO 0);
SIGNAL \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|locked_wire\ : std_logic_vector(0 DOWNTO 0);
SIGNAL \TheRxFsk|ALT_INV_Add2~37_sumout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Add2~33_sumout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Add2~29_sumout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Add2~25_sumout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Add2~21_sumout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Add2~17_sumout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Add2~13_sumout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Add2~9_sumout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Add2~5_sumout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Add2~1_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Add4~17_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Sum[-2]~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_DdryDelayed\ : std_logic_vector(0 DOWNTO 0);
SIGNAL \TheRxFsk|Lowpass|ALT_INV_DdryDelayed[-1]~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_DdryDelayed[-2]~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_DdryDelayed[-3]~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_DdryDelayed[-4]~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_DdryDelayed[-5]~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_DdryDelayed[-6]~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_DdryDelayed[-7]~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_DdryDelayed[-8]~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_DdryDelayed[-9]~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_DdryDelayed[-10]~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_DdryDelayed[-11]~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_DdryDelayed[-12]~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_DdryDelayed[-13]~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_DdryDelayed[-14]~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_DdryDelayed[-15]~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a1\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a2\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a3\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a4\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a5\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a6\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a7\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a8\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a9\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a10\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a11\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a12\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a13\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a14\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a15\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a0~portbdataout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Add4~13_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Sum[-1]~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Mult0~39\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Mult0~38\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Mult0~37\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Mult0~36\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Mult0~35\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Mult0~34\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Mult0~33\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Mult0~32\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Mult0~31\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Mult0~30\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Mult0~29\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Mult0~28\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Mult0~27\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Mult0~26\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Mult0~25\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Mult0~24\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Mult0~23\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Mult0~22\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Mult0~21\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Mult0~20\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Mult0~19\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Mult0~18\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Mult0~17\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Mult0~16\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Mult0~15\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Mult0~14\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Mult0~13\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Mult0~12\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Mult0~11\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Mult0~10\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Mult0~9\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Mult0~8_resulta\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Add2~25_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Add2~21_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Add2~13_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Add2~9_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Add2~5_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Add2~1_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Add4~9_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Add3~1_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Add4~5_sumout\ : std_logic;
SIGNAL \GenClks|ALT_INV_Add0~29_sumout\ : std_logic;
SIGNAL \GenClks|ALT_INV_Add0~13_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Add4~1_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Sum\ : std_logic_vector(0 DOWNTO 0);
SIGNAL \ConfigureCodec|ALT_INV_R.AddrCtr\ : std_logic_vector(6 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.EnableSumUp~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.SelSumUp~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_R.EnableSumUp~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_R.SelSumUp~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_R.EnableSumUp~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_R.SelSumUp~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_R.EnableSumUp~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_R.SelSumUp~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_MultResult[-4]~3_combout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Mux1~0_combout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Mux17~0_combout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Mux2~0_combout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Mux18~0_combout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Mux3~0_combout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Mux19~0_combout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Mux4~0_combout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Mux20~0_combout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Mux5~0_combout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Mux21~0_combout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Mux6~0_combout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Mux22~0_combout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Mux7~0_combout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Mux23~0_combout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Mux8~0_combout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Mux24~0_combout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Mux9~0_combout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Mux25~0_combout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Mux10~0_combout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Mux26~0_combout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Mux11~0_combout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Mux27~0_combout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Mux12~0_combout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Mux28~0_combout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Mux13~0_combout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Mux29~0_combout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Mux14~0_combout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Mux30~0_combout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Mux15~0_combout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Mux31~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:11:Bandpass0|ALT_INV_R.SumState.Idle~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_MultResult[-3]~2_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Equal0~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Equal2~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.AddressState~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:11:Bandpass0|ALT_INV_R.SumState.SumEnable~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_MultResult[-2]~1_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressSample\ : std_logic_vector(6 DOWNTO 0);
SIGNAL \TheRxFsk|Lowpass|ALT_INV_R.WriteAddress\ : std_logic_vector(6 DOWNTO 0);
SIGNAL \TheRxFsk|Lowpass|ALT_INV_CoefMemory~7_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_CoefMemory~5_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_CoefMemory~4_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_CoefMemory~2_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_CoefMemory~1_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:11:Bandpass1|ALT_INV_Equal1~1_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.ReadAddressCoef\ : std_logic_vector(8 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:11:Bandpass1|ALT_INV_Equal1~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:11:Bandpass0|ALT_INV_R.SumState.SumSelect~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_MultResult[-1]~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_R.FirstSample~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_R.AddressState~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:11:Bandpass0|ALT_INV_R.SumState.SumWait2~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:11:Bandpass0|ALT_INV_R.SumState.SumValid~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Equal1~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\ : std_logic_vector(6 DOWNTO 0);
SIGNAL \TheRxFsk|Lowpass|ALT_INV_R.SumState.SumSelect~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_CoefMemory~0_combout\ : std_logic;
SIGNAL \ConfigureCodec|ALT_INV_Selector13~2_combout\ : std_logic;
SIGNAL \ConfigureCodec|ALT_INV_Selector12~1_combout\ : std_logic;
SIGNAL \ConfigureCodec|ALT_INV_Selector12~0_combout\ : std_logic;
SIGNAL \ConfigureCodec|ALT_INV_Selector11~2_combout\ : std_logic;
SIGNAL \ConfigureCodec|ALT_INV_NextR~10_combout\ : std_logic;
SIGNAL \ConfigureCodec|ALT_INV_Mux8~0_combout\ : std_logic;
SIGNAL \ConfigureCodec|ALT_INV_Selector11~1_combout\ : std_logic;
SIGNAL \ConfigureCodec|ALT_INV_Selector11~0_combout\ : std_logic;
SIGNAL \ConfigureCodec|ALT_INV_Selector10~1_combout\ : std_logic;
SIGNAL \ConfigureCodec|ALT_INV_Selector5~0_combout\ : std_logic;
SIGNAL \ConfigureCodec|ALT_INV_Selector10~0_combout\ : std_logic;
SIGNAL \ConfigureCodec|ALT_INV_Selector13~1_combout\ : std_logic;
SIGNAL \ConfigureCodec|ALT_INV_Selector1~0_combout\ : std_logic;
SIGNAL \ConfigureCodec|ALT_INV_Selector15~2_combout\ : std_logic;
SIGNAL \ConfigureCodec|ALT_INV_Selector15~1_combout\ : std_logic;
SIGNAL \ConfigureCodec|ALT_INV_R.FrameState.Start~q\ : std_logic;
SIGNAL \ConfigureCodec|ALT_INV_Selector15~0_combout\ : std_logic;
SIGNAL \ConfigureCodec|ALT_INV_R.FrameState.Address~q\ : std_logic;
SIGNAL \ConfigureCodec|ALT_INV_Mux9~4_combout\ : std_logic;
SIGNAL \ConfigureCodec|ALT_INV_Mux9~3_combout\ : std_logic;
SIGNAL \ConfigureCodec|ALT_INV_R.Data\ : std_logic_vector(15 DOWNTO 0);
SIGNAL \ConfigureCodec|ALT_INV_Mux9~2_combout\ : std_logic;
SIGNAL \ConfigureCodec|ALT_INV_Mux9~1_combout\ : std_logic;
SIGNAL \ConfigureCodec|ALT_INV_Mux9~0_combout\ : std_logic;
SIGNAL \TheI2sToPar|ALT_INV_LrcDlyd~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_R.SumState.Idle~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:11:Bandpass0|ALT_INV_R.ValWet~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_R.SumState.SumEnable~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed\ : std_logic_vector(0 DOWNTO 0);
SIGNAL \ConfigureCodec|ALT_INV_R.FrameState.Data1~q\ : std_logic;
SIGNAL \ConfigureCodec|ALT_INV_NextR~9_combout\ : std_logic;
SIGNAL \ConfigureCodec|ALT_INV_R.FrameState.RWBit~q\ : std_logic;
SIGNAL \ConfigureCodec|ALT_INV_NextR~8_combout\ : std_logic;
SIGNAL \ConfigureCodec|ALT_INV_R.BitCtr\ : std_logic_vector(3 DOWNTO 0);
SIGNAL \ConfigureCodec|ALT_INV_R.FrameState.Data2~q\ : std_logic;
SIGNAL \ConfigureCodec|ALT_INV_R.Sdin~q\ : std_logic;
SIGNAL \TheI2sToPar|ALT_INV_Decoder0~4_combout\ : std_logic;
SIGNAL \TheI2sToPar|ALT_INV_D[14]~7_combout\ : std_logic;
SIGNAL \TheI2sToPar|ALT_INV_Decoder0~3_combout\ : std_logic;
SIGNAL \TheI2sToPar|ALT_INV_Decoder0~2_combout\ : std_logic;
SIGNAL \TheI2sToPar|ALT_INV_Decoder0~1_combout\ : std_logic;
SIGNAL \TheI2sToPar|ALT_INV_Equal0~2_combout\ : std_logic;
SIGNAL \TheI2sToPar|ALT_INV_Equal0~1_combout\ : std_logic;
SIGNAL \TheI2sToPar|ALT_INV_BclkRiseEdge~combout\ : std_logic;
SIGNAL \TheI2sToPar|ALT_INV_Equal0~0_combout\ : std_logic;
SIGNAL \TheI2sToPar|ALT_INV_AudioBitCtr\ : std_logic_vector(4 DOWNTO 0);
SIGNAL \TheI2sToPar|ALT_INV_Decoder0~0_combout\ : std_logic;
SIGNAL \TheI2sToPar|ALT_INV_State~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_R.EnableSumUp~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_R.SelSumUp~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_R.SumState.SumWait2~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_R.SumState.SumValid~q\ : std_logic;
SIGNAL \ConfigureCodec|ALT_INV_NextStateAndOutput:vSclkFalling~0_combout\ : std_logic;
SIGNAL \ConfigureCodec|ALT_INV_Selector13~0_combout\ : std_logic;
SIGNAL \ConfigureCodec|ALT_INV_R.FrameState.Ack2~q\ : std_logic;
SIGNAL \ConfigureCodec|ALT_INV_R.FrameState.Ack1~q\ : std_logic;
SIGNAL \ConfigureCodec|ALT_INV_R.FrameState.Ack3~q\ : std_logic;
SIGNAL \ConfigureCodec|ALT_INV_R.Activity~0_combout\ : std_logic;
SIGNAL \ConfigureCodec|ALT_INV_Selector16~0_combout\ : std_logic;
SIGNAL \GenStrobeI2C|ALT_INV_ClkCounter\ : std_logic_vector(5 DOWNTO 0);
SIGNAL \GenClks|ALT_INV_Equal0~0_combout\ : std_logic;
SIGNAL \GenClks|ALT_INV_BitCounter\ : std_logic_vector(7 DOWNTO 0);
SIGNAL \GenClks|ALT_INV_ADClrc~0_combout\ : std_logic;
SIGNAL \TheParToI2s|ALT_INV_NextState~6_combout\ : std_logic;
SIGNAL \TheParToI2s|ALT_INV_Selector9~0_combout\ : std_logic;
SIGNAL \TheParToI2s|ALT_INV_Selector7~0_combout\ : std_logic;
SIGNAL \TheParToI2s|ALT_INV_Add0~0_combout\ : std_logic;
SIGNAL \TheI2sToPar|ALT_INV_D\ : std_logic_vector(15 DOWNTO 0);
SIGNAL \TheParToI2s|ALT_INV_Selector8~0_combout\ : std_logic;
SIGNAL \TheParToI2s|ALT_INV_NextBclkCtr~1_combout\ : std_logic;
SIGNAL \TheParToI2s|ALT_INV_Selector6~1_combout\ : std_logic;
SIGNAL \TheParToI2s|ALT_INV_NextBclkCtr~0_combout\ : std_logic;
SIGNAL \TheParToI2s|ALT_INV_State.SyncingToBclk~q\ : std_logic;
SIGNAL \TheParToI2s|ALT_INV_State.WaitingValL~q\ : std_logic;
SIGNAL \TheParToI2s|ALT_INV_Selector6~0_combout\ : std_logic;
SIGNAL \TheI2sToPar|ALT_INV_BclkDlyd~q\ : std_logic;
SIGNAL \TheParToI2s|ALT_INV_State.FirstBitEmptyR~q\ : std_logic;
SIGNAL \TheI2sToPar|ALT_INV_ValL~q\ : std_logic;
SIGNAL \GenClks|ALT_INV_ClkCounter\ : std_logic_vector(0 DOWNTO 0);
SIGNAL \TheRxFsk|Lowpass|ALT_INV_R.ValWet~q\ : std_logic;
SIGNAL \ConfigureCodec|ALT_INV_R.AddrCtr[6]~1_combout\ : std_logic;
SIGNAL \ConfigureCodec|ALT_INV_R.FrameState.Stop~q\ : std_logic;
SIGNAL \ConfigureCodec|ALT_INV_R.AckError~q\ : std_logic;
SIGNAL \ConfigureCodec|ALT_INV_R.Sclk~q\ : std_logic;
SIGNAL \ConfigureCodec|ALT_INV_Equal0~1_combout\ : std_logic;
SIGNAL \ConfigureCodec|ALT_INV_R.AddrCtr[6]~0_combout\ : std_logic;
SIGNAL \ConfigureCodec|ALT_INV_R.FrameState.Idle~q\ : std_logic;
SIGNAL \ConfigureCodec|ALT_INV_R.Activity~q\ : std_logic;
SIGNAL \ConfigureCodec|ALT_INV_Equal0~0_combout\ : std_logic;
SIGNAL ALT_INV_WaitCtr : std_logic_vector(1 DOWNTO 0);
SIGNAL \GenStrobeI2C|ALT_INV_oStrobe~q\ : std_logic;
SIGNAL \TheParToI2s|ALT_INV_oLrc~0_combout\ : std_logic;
SIGNAL \TheParToI2s|ALT_INV_State.FirstBitEmptyL~q\ : std_logic;
SIGNAL \GenClks|ALT_INV_ADClrc~q\ : std_logic;
SIGNAL \TheParToI2s|ALT_INV_Selector10~0_combout\ : std_logic;
SIGNAL \TheParToI2s|ALT_INV_State.SendingR~q\ : std_logic;
SIGNAL \TheParToI2s|ALT_INV_State.SendingL~q\ : std_logic;
SIGNAL \TheParToI2s|ALT_INV_BclkCtr\ : std_logic_vector(3 DOWNTO 0);
SIGNAL \TheParToI2s|ALT_INV_Mux1~3_combout\ : std_logic;
SIGNAL \TheParToI2s|ALT_INV_LastValidDL\ : std_logic_vector(15 DOWNTO 0);
SIGNAL \TheParToI2s|ALT_INV_Mux1~2_combout\ : std_logic;
SIGNAL \TheParToI2s|ALT_INV_Mux1~1_combout\ : std_logic;
SIGNAL \TheParToI2s|ALT_INV_Mux1~0_combout\ : std_logic;
SIGNAL \GenClks|ALT_INV_BMclk~q\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_oD~q\ : std_logic;
SIGNAL \ConfigureCodec|ALT_INV_R.Configured~q\ : std_logic;
SIGNAL \ALT_INV_Start~q\ : std_logic;
SIGNAL \SyncSwitchInput|ALT_INV_Metastable\ : std_logic_vector(1 DOWNTO 1);
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Sum[-15]~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Sum[-14]~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Add4~61_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Sum[-13]~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Add4~57_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Sum[-12]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add0~33_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add0~5_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add1~33_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Add4~53_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Sum[-11]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.WriteAddress\ : std_logic_vector(8 DOWNTO 0);
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Add4~49_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Sum[-10]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a13\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a14\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a15\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a1\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a2\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a3\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a4\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a5\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a6\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a7\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a8\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a9\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a12~portbdataout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a10\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a8\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a9\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a11\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a10\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a11\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a12\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a13\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a14\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a15\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a0~portbdataout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a5\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a6\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a7\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a8\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a9\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a10\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a11\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a12\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a13\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a14\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a0\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a1\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a2\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a3\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a4\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a5\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a6\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a7\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a15\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a1\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a2\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a3\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a0\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a1\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a2\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a3\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a4\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a5\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a6\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a7\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a8\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a9\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a4~portbdataout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a10\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a11\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a12\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a13\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a14\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a15\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a0~portbdataout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Add4~45_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Sum[-9]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~39\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~38\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~37\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~36\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~35\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~34\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~33\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~32\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~31\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~30\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~29\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~28\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~27\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~26\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~25\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~24\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~23\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~22\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~21\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~20\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~19\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~18\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~17\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~16\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~15\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~14\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~13\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~12\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~11\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~10\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~9\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~8_resulta\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~39\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~38\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~37\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~36\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~35\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~34\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~33\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~32\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~31\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~30\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~29\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~28\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~27\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~26\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~25\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~24\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~23\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~22\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~21\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~20\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~19\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~18\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~17\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~16\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~15\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~14\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~13\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~12\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~11\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~10\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~9\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~8_resulta\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~39\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~38\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~37\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~36\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~35\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~34\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~33\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~32\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~31\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~30\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~29\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~28\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~27\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~26\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~25\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~24\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~23\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~22\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~21\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~20\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~19\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~18\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~17\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~16\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~15\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~14\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~13\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~12\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~11\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~10\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~9\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~8_resulta\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~39\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~38\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~37\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~36\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~35\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~34\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~33\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~32\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~31\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~30\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~29\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~28\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~27\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~26\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~25\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~24\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~23\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~22\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~21\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~20\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~19\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~18\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~17\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~16\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~15\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~14\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~13\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~12\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~11\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~10\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~9\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~8_resulta\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Add4~41_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Sum[-8]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add3~1_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add3~1_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add3~1_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add3~1_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Add4~37_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Sum[-7]~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Add4~33_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Sum[-6]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~65_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~65_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~65_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~65_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~61_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~61_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~61_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~61_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~57_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~57_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~57_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~57_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~53_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~53_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~53_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~53_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~49_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~49_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~49_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~49_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~45_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~45_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~45_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~45_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~41_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~41_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~41_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~41_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~37_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~37_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~37_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~37_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~33_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~33_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~33_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~33_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~29_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~29_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~29_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~29_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~25_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~25_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~25_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~25_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~21_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~21_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~21_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~21_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~17_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~17_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~17_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~17_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~13_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~13_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~13_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~13_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~5_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~5_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~1_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~1_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~5_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~5_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~1_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~1_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Add4~29_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Sum[-5]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-1]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-1]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-1]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-1]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-2]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-2]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-2]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-2]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-3]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-3]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-3]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-3]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-4]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-4]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-4]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-4]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-5]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-5]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-5]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-5]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-6]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-6]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-6]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-6]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-7]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-7]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-7]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-7]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-8]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-8]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-8]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-8]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-9]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-9]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-9]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-9]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-10]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-10]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-10]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-10]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-11]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-11]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-11]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-11]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-12]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-12]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-12]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-12]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-13]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-13]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-13]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-13]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-14]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-14]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-14]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-14]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-15]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-15]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum\ : std_logic_vector(0 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum\ : std_logic_vector(0 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-15]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-15]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum\ : std_logic_vector(0 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum\ : std_logic_vector(0 DOWNTO 0);
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Add4~25_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Sum[-4]~q\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Add0~61_sumout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Add1~61_sumout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Add0~57_sumout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Add1~57_sumout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Add0~53_sumout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Add1~53_sumout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Add0~49_sumout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Add1~49_sumout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Add0~45_sumout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Add1~45_sumout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Add0~41_sumout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Add1~41_sumout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Add0~37_sumout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Add1~37_sumout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Add0~33_sumout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Add1~33_sumout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Add0~29_sumout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Add1~29_sumout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Add0~25_sumout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Add1~25_sumout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Add0~21_sumout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Add1~21_sumout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Add0~17_sumout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Add1~17_sumout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Add0~13_sumout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Add1~13_sumout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Add0~9_sumout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Add1~9_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Add0~25_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Add0~13_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Add0~5_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Add1~25_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Add1~21_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Add1~17_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Add1~13_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Add1~9_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Add1~5_sumout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Add0~5_sumout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Add1~5_sumout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Add0~1_sumout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Add1~1_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_Add2~29_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_Add2~25_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_Add2~21_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_Add2~17_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_Add2~13_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_Add2~9_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_Add2~5_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_Add2~1_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Add4~21_sumout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_Sum[-3]~q\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Add2~65_sumout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Add2~61_sumout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Add2~57_sumout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Add2~53_sumout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Add2~49_sumout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Add2~45_sumout\ : std_logic;
SIGNAL \TheRxFsk|ALT_INV_Add2~41_sumout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[0]~DUPLICATE_q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_R.SumState.Idle~DUPLICATE_q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_R.SumState.SumEnable~DUPLICATE_q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressSample[0]~DUPLICATE_q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_R.WriteAddress[1]~DUPLICATE_q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.ReadAddressCoef[0]~DUPLICATE_q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.ReadAddressCoef[1]~DUPLICATE_q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.ReadAddressCoef[2]~DUPLICATE_q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.ReadAddressCoef[4]~DUPLICATE_q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.ReadAddressCoef[5]~DUPLICATE_q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.ReadAddressCoef[6]~DUPLICATE_q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.ReadAddressCoef[7]~DUPLICATE_q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef[6]~DUPLICATE_q\ : std_logic;
SIGNAL \ConfigureCodec|ALT_INV_R.FrameState.Data1~DUPLICATE_q\ : std_logic;
SIGNAL \ConfigureCodec|ALT_INV_R.BitCtr[0]~DUPLICATE_q\ : std_logic;
SIGNAL \ConfigureCodec|ALT_INV_R.BitCtr[3]~DUPLICATE_q\ : std_logic;
SIGNAL \ConfigureCodec|ALT_INV_R.FrameState.Data2~DUPLICATE_q\ : std_logic;
SIGNAL \TheI2sToPar|ALT_INV_AudioBitCtr[1]~DUPLICATE_q\ : std_logic;
SIGNAL \TheI2sToPar|ALT_INV_AudioBitCtr[2]~DUPLICATE_q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_R.SumState.SumWait2~DUPLICATE_q\ : std_logic;
SIGNAL \ConfigureCodec|ALT_INV_R.FrameState.Ack1~DUPLICATE_q\ : std_logic;
SIGNAL \GenStrobeI2C|ALT_INV_ClkCounter[0]~DUPLICATE_q\ : std_logic;
SIGNAL \GenStrobeI2C|ALT_INV_ClkCounter[1]~DUPLICATE_q\ : std_logic;
SIGNAL \GenClks|ALT_INV_BitCounter[1]~DUPLICATE_q\ : std_logic;
SIGNAL \TheParToI2s|ALT_INV_State.SyncingToBclk~DUPLICATE_q\ : std_logic;
SIGNAL \ConfigureCodec|ALT_INV_R.FrameState.Idle~DUPLICATE_q\ : std_logic;
SIGNAL \ALT_INV_WaitCtr[0]~DUPLICATE_q\ : std_logic;
SIGNAL \TheParToI2s|ALT_INV_BclkCtr[2]~DUPLICATE_q\ : std_logic;
SIGNAL \TheParToI2s|ALT_INV_BclkCtr[3]~DUPLICATE_q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-2]~DUPLICATE_q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-3]~DUPLICATE_q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-3]~DUPLICATE_q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-4]~DUPLICATE_q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-7]~DUPLICATE_q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-8]~DUPLICATE_q\ : std_logic;
SIGNAL \ConfigureCodec|ALT_INV_R.AddrCtr[1]~DUPLICATE_q\ : std_logic;
SIGNAL \ConfigureCodec|ALT_INV_R.AddrCtr[2]~DUPLICATE_q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-14]_OTERM179\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-14]_OTERM177\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-14]_OTERM175\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-13]_OTERM173\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-13]_OTERM171\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-13]_OTERM169\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-12]_OTERM167\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-12]_OTERM165\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-12]_OTERM163\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-11]_OTERM161\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-11]_OTERM159\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-11]_OTERM157\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-10]_OTERM155\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-10]_OTERM153\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-10]_OTERM151\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-9]_OTERM149\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-9]_OTERM147\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-9]_OTERM145\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-8]_OTERM143\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-8]_OTERM141\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-8]_OTERM139\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-7]_OTERM137\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-7]_OTERM135\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-7]_OTERM133\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-6]_OTERM131\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-6]_OTERM129\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-6]_OTERM127\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-5]_OTERM125\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-5]_OTERM123\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-5]_OTERM121\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-4]_OTERM119\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-4]_OTERM117\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-4]_OTERM115\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-3]_OTERM113\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-3]_OTERM111\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-3]_OTERM109\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-2]_OTERM107\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-2]_OTERM105\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-2]_OTERM103\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-1]_OTERM101\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-1]_OTERM99\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-1]_OTERM97\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-14]_OTERM95\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-14]_OTERM93\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-13]_OTERM91\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-13]_OTERM89\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM87\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM85\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM83\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM81\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM79\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM77\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM75\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM73\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM71\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM69\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM67\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM65\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-12]_OTERM63\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-12]_OTERM61\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-11]_OTERM59\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-11]_OTERM57\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-10]_OTERM55\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-9]_OTERM53\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-9]_OTERM51\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-10]_OTERM49\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-8]_OTERM47\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-8]_OTERM45\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-7]_OTERM43\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-7]_OTERM41\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-6]_OTERM39\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-6]_OTERM37\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-5]_OTERM35\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-5]_OTERM33\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-4]_OTERM31\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-4]_OTERM29\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-3]_OTERM27\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-3]_OTERM25\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-2]_OTERM23\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-2]_OTERM21\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-1]_OTERM19\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-1]_OTERM17\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM15\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM13\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM11\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM9\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM7\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM5\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM3\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM1\ : std_logic;
SIGNAL \ALT_INV_iADCdat~input_o\ : std_logic;
SIGNAL \ALT_INV_inResetAsync~input_o\ : std_logic;
SIGNAL \ALT_INV_ioI2cSdin~input_o\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_CoefMemory~34_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_CoefMemory~33_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_CoefMemory~31_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_CoefMemory~30_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_CoefMemory~28_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_CoefMemory~27_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_CoefMemory~25_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_CoefMemory~24_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_CoefMemory~22_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_CoefMemory~21_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_CoefMemory~19_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_CoefMemory~18_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_CoefMemory~16_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_CoefMemory~15_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_CoefMemory~13_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_CoefMemory~12_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_CoefMemory~10_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_CoefMemory~9_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_vAdd~2_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_vAdd~1_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_vAdd~2_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_vAdd~1_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_vAdd~2_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_vAdd~1_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_vAdd~2_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_vAdd~1_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_vAdd~2_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_vAdd~1_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_vAdd~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_MultResult[-15]~14_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_MultResult[-14]~13_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_MultResult[-13]~12_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_MultResult[-12]~11_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_MultResult[-11]~10_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Equal0~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Equal2~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_MultResult[-10]~9_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.ReadAddressSample\ : std_logic_vector(8 DOWNTO 0);
SIGNAL \TheRxFsk|Lowpass|ALT_INV_MultResult[-9]~8_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed\ : std_logic_vector(0 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-1]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-2]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-3]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-4]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-5]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-6]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-7]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-8]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-9]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-10]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-11]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-12]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-13]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-14]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-15]~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_MultResult[-8]~7_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_vAdd~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_vAdd~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.SumState.SumSelect~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_R.SumState.SumSelect~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_vAdd~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_vAdd~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_R.SumState.SumSelect~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_R.SumState.SumSelect~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_MultResult[-7]~6_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResult[-1]~14_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResult[-1]~14_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResult[-1]~14_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResult[-1]~14_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResult[-2]~13_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResult[-2]~13_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResult[-2]~13_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResult[-2]~13_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResult[-3]~12_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResult[-3]~12_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResult[-3]~12_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResult[-3]~12_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResult[-4]~11_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResult[-4]~11_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResult[-4]~11_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResult[-4]~11_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResult[-5]~10_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResult[-5]~10_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResult[-5]~10_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResult[-5]~10_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResult[-6]~9_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResult[-6]~9_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResult[-6]~9_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResult[-6]~9_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResult[-7]~8_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResult[-7]~8_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResult[-7]~8_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResult[-7]~8_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResult[-8]~7_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResult[-8]~7_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResult[-8]~7_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResult[-8]~7_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResult[-9]~6_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResult[-9]~6_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResult[-9]~6_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResult[-9]~6_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResult[-10]~5_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResult[-10]~5_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResult[-10]~5_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResult[-10]~5_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResult[-11]~4_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResult[-11]~4_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResult[-11]~4_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResult[-11]~4_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResult[-12]~3_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResult[-12]~3_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResult[-12]~3_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResult[-12]~3_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResult[-13]~2_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResult[-13]~2_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResult[-13]~2_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResult[-13]~2_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResult[-14]~1_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResult[-14]~1_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResult[-14]~1_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResult[-14]~1_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResult[-15]~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResult[-15]~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.SumState.SumValid~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_R.SumState.SumValid~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResult[-15]~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResult[-15]~0_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_R.SumState.SumValid~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_R.SumState.SumValid~q\ : std_logic;
SIGNAL \TheRxFsk|Lowpass|ALT_INV_MultResult[-6]~5_combout\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.SumState.Idle~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.SumState.SumEnable~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.SumState.SumWait2~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed\ : std_logic_vector(0 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_R.SumState.Idle~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_R.SumState.SumEnable~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_R.SumState.SumWait2~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed\ : std_logic_vector(0 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_R.SumState.Idle~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_R.SumState.SumEnable~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_R.SumState.SumWait2~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed\ : std_logic_vector(0 DOWNTO 0);
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_R.SumState.Idle~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_R.SumState.SumEnable~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_R.SumState.SumWait2~q\ : std_logic;
SIGNAL \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed\ : std_logic_vector(0 DOWNTO 0);
SIGNAL \TheRxFsk|Lowpass|ALT_INV_MultResult[-5]~4_combout\ : std_logic;

BEGIN

ww_iClk <= iClk;
ww_inResetAsync <= inResetAsync;
ww_iSwitch <= IEEE.STD_LOGIC_1164.TO_STDLOGICVECTOR(iSwitch);
ww_inButton <= IEEE.STD_LOGIC_1164.TO_STDLOGICVECTOR(inButton);
oSEG0 <= IEEE.STD_LOGIC_1164.TO_STDULOGICVECTOR(ww_oSEG0);
oSEG1 <= IEEE.STD_LOGIC_1164.TO_STDULOGICVECTOR(ww_oSEG1);
oSEG2 <= IEEE.STD_LOGIC_1164.TO_STDULOGICVECTOR(ww_oSEG2);
oSEG3 <= IEEE.STD_LOGIC_1164.TO_STDULOGICVECTOR(ww_oSEG3);
oSEG4 <= IEEE.STD_LOGIC_1164.TO_STDULOGICVECTOR(ww_oSEG4);
oSEG5 <= IEEE.STD_LOGIC_1164.TO_STDULOGICVECTOR(ww_oSEG5);
oLed <= IEEE.STD_LOGIC_1164.TO_STDULOGICVECTOR(ww_oLed);
oI2cSclk <= ww_oI2cSclk;
oMclk <= ww_oMclk;
oBclk <= ww_oBclk;
ww_iADCdat <= iADCdat;
oDACdat <= ww_oDACdat;
oADClrc <= ww_oADClrc;
oDAClrc <= ww_oDAClrc;
ww_devoe <= devoe;
ww_devclrn <= devclrn;
ww_devpor <= devpor;

\TheRxFsk|Lowpass|Mult0~8_ACLR_bus\ <= (gnd & gnd);

\TheRxFsk|Lowpass|Mult0~8_CLK_bus\ <= (gnd & gnd & \iClk~inputCLKENA0_outclk\);

\TheRxFsk|Lowpass|Mult0~8_ENA_bus\ <= (vcc & vcc & vcc);

\TheRxFsk|Lowpass|Mult0~8_AX_bus\ <= (\TheRxFsk|Lowpass|CoefMemory~8_combout\ & \TheRxFsk|Lowpass|CoefMemory~8_combout\ & \TheRxFsk|Lowpass|CoefMemory~8_combout\ & \TheRxFsk|Lowpass|CoefMemory~8_combout\ & \TheRxFsk|Lowpass|CoefMemory~8_combout\ & 
\TheRxFsk|Lowpass|CoefMemory~8_combout\ & \TheRxFsk|Lowpass|CoefMemory~8_combout\ & \TheRxFsk|Lowpass|CoefMemory~6_combout\ & \TheRxFsk|Lowpass|CoefMemory~3_combout\ & \TheRxFsk|Lowpass|CoefMemory~11_combout\ & \TheRxFsk|Lowpass|CoefMemory~14_combout\ & 
\TheRxFsk|Lowpass|CoefMemory~17_combout\ & \TheRxFsk|Lowpass|CoefMemory~20_combout\ & \TheRxFsk|Lowpass|CoefMemory~23_combout\ & \TheRxFsk|Lowpass|CoefMemory~26_combout\ & \TheRxFsk|Lowpass|CoefMemory~29_combout\ & \TheRxFsk|Lowpass|CoefMemory~32_combout\
& \TheRxFsk|Lowpass|CoefMemory~35_combout\);

\TheRxFsk|Lowpass|Mult0~8_AY_bus\ <= (\TheRxFsk|Lowpass|Sample[0]~15_combout\ & \TheRxFsk|Lowpass|Sample[0]~15_combout\ & \TheRxFsk|Lowpass|Sample[0]~15_combout\ & \TheRxFsk|Lowpass|Sample[0]~15_combout\ & \TheRxFsk|Lowpass|Sample[-1]~14_combout\ & 
\TheRxFsk|Lowpass|Sample[-2]~13_combout\ & \TheRxFsk|Lowpass|Sample[-3]~12_combout\ & \TheRxFsk|Lowpass|Sample[-4]~11_combout\ & \TheRxFsk|Lowpass|Sample[-5]~10_combout\ & \TheRxFsk|Lowpass|Sample[-6]~9_combout\ & \TheRxFsk|Lowpass|Sample[-7]~8_combout\
& \TheRxFsk|Lowpass|Sample[-8]~7_combout\ & \TheRxFsk|Lowpass|Sample[-9]~6_combout\ & \TheRxFsk|Lowpass|Sample[-10]~5_combout\ & \TheRxFsk|Lowpass|Sample[-11]~4_combout\ & \TheRxFsk|Lowpass|Sample[-12]~3_combout\ & \TheRxFsk|Lowpass|Sample[-13]~2_combout\
& \TheRxFsk|Lowpass|Sample[-14]~1_combout\ & \TheRxFsk|Lowpass|Sample[-15]~0_combout\);

\TheRxFsk|Lowpass|Mult0~8_resulta\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(0);
\TheRxFsk|Lowpass|Mult0~9\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(1);
\TheRxFsk|Lowpass|Mult0~10\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(2);
\TheRxFsk|Lowpass|Mult0~11\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(3);
\TheRxFsk|Lowpass|Mult0~12\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(4);
\TheRxFsk|Lowpass|Mult0~13\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(5);
\TheRxFsk|Lowpass|Mult0~14\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(6);
\TheRxFsk|Lowpass|Mult0~15\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(7);
\TheRxFsk|Lowpass|Mult0~16\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(8);
\TheRxFsk|Lowpass|Mult0~17\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(9);
\TheRxFsk|Lowpass|Mult0~18\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(10);
\TheRxFsk|Lowpass|Mult0~19\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(11);
\TheRxFsk|Lowpass|Mult0~20\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(12);
\TheRxFsk|Lowpass|Mult0~21\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(13);
\TheRxFsk|Lowpass|Mult0~22\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(14);
\TheRxFsk|Lowpass|Mult0~23\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(15);
\TheRxFsk|Lowpass|Mult0~24\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(16);
\TheRxFsk|Lowpass|Mult0~25\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(17);
\TheRxFsk|Lowpass|Mult0~26\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(18);
\TheRxFsk|Lowpass|Mult0~27\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(19);
\TheRxFsk|Lowpass|Mult0~28\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(20);
\TheRxFsk|Lowpass|Mult0~29\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(21);
\TheRxFsk|Lowpass|Mult0~30\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(22);
\TheRxFsk|Lowpass|Mult0~31\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(23);
\TheRxFsk|Lowpass|Mult0~32\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(24);
\TheRxFsk|Lowpass|Mult0~33\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(25);
\TheRxFsk|Lowpass|Mult0~34\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(26);
\TheRxFsk|Lowpass|Mult0~35\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(27);
\TheRxFsk|Lowpass|Mult0~36\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(28);
\TheRxFsk|Lowpass|Mult0~37\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(29);
\TheRxFsk|Lowpass|Mult0~38\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(30);
\TheRxFsk|Lowpass|Mult0~39\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(31);
\TheRxFsk|Lowpass|Mult0~40\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(32);
\TheRxFsk|Lowpass|Mult0~41\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(33);
\TheRxFsk|Lowpass|Mult0~42\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(34);
\TheRxFsk|Lowpass|Mult0~43\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(35);
\TheRxFsk|Lowpass|Mult0~44\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(36);
\TheRxFsk|Lowpass|Mult0~45\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(37);
\TheRxFsk|Lowpass|Mult0~46\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(38);
\TheRxFsk|Lowpass|Mult0~47\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(39);
\TheRxFsk|Lowpass|Mult0~48\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(40);
\TheRxFsk|Lowpass|Mult0~49\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(41);
\TheRxFsk|Lowpass|Mult0~50\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(42);
\TheRxFsk|Lowpass|Mult0~51\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(43);
\TheRxFsk|Lowpass|Mult0~52\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(44);
\TheRxFsk|Lowpass|Mult0~53\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(45);
\TheRxFsk|Lowpass|Mult0~54\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(46);
\TheRxFsk|Lowpass|Mult0~55\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(47);
\TheRxFsk|Lowpass|Mult0~56\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(48);
\TheRxFsk|Lowpass|Mult0~57\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(49);
\TheRxFsk|Lowpass|Mult0~58\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(50);
\TheRxFsk|Lowpass|Mult0~59\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(51);
\TheRxFsk|Lowpass|Mult0~60\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(52);
\TheRxFsk|Lowpass|Mult0~61\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(53);
\TheRxFsk|Lowpass|Mult0~62\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(54);
\TheRxFsk|Lowpass|Mult0~63\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(55);
\TheRxFsk|Lowpass|Mult0~64\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(56);
\TheRxFsk|Lowpass|Mult0~65\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(57);
\TheRxFsk|Lowpass|Mult0~66\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(58);
\TheRxFsk|Lowpass|Mult0~67\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(59);
\TheRxFsk|Lowpass|Mult0~68\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(60);
\TheRxFsk|Lowpass|Mult0~69\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(61);
\TheRxFsk|Lowpass|Mult0~70\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(62);
\TheRxFsk|Lowpass|Mult0~71\ <= \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\(63);

\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTADATAIN_bus\ <= (gnd & gnd & gnd & gnd & gnd & gnd & gnd & gnd & gnd & gnd & gnd & gnd & gnd & gnd & gnd & gnd & gnd & gnd & gnd & gnd & gnd & gnd & gnd & gnd & \TheRxFsk|Add2~5_sumout\
& \TheRxFsk|Substracted[-1]~14_combout\ & \TheRxFsk|Substracted[-2]~13_combout\ & \TheRxFsk|Substracted[-3]~12_combout\ & \TheRxFsk|Substracted[-4]~11_combout\ & \TheRxFsk|Substracted[-5]~10_combout\ & \TheRxFsk|Substracted[-6]~9_combout\ & 
\TheRxFsk|Substracted[-7]~8_combout\ & \TheRxFsk|Substracted[-8]~7_combout\ & \TheRxFsk|Substracted[-9]~6_combout\ & \TheRxFsk|Substracted[-10]~5_combout\ & \TheRxFsk|Substracted[-11]~4_combout\ & \TheRxFsk|Substracted[-12]~3_combout\ & 
\TheRxFsk|Substracted[-13]~2_combout\ & \TheRxFsk|Substracted[-14]~1_combout\ & \TheRxFsk|Substracted[-15]~0_combout\);

\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTAADDR_bus\ <= (\TheRxFsk|Lowpass|R.WriteAddress[6]~_wirecell_combout\ & \TheRxFsk|Lowpass|R.WriteAddress\(5) & \TheRxFsk|Lowpass|R.WriteAddress\(4) & 
\TheRxFsk|Lowpass|R.WriteAddress[3]~_wirecell_combout\ & \TheRxFsk|Lowpass|R.WriteAddress\(2) & \TheRxFsk|Lowpass|R.WriteAddress[1]~_wirecell_combout\ & \TheRxFsk|Lowpass|R.WriteAddress[0]~DUPLICATE_q\);

\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBADDR_bus\ <= (\TheRxFsk|Lowpass|R.ReadAddressSample\(6) & \TheRxFsk|Lowpass|R.ReadAddressSample\(5) & \TheRxFsk|Lowpass|R.ReadAddressSample\(4) & 
\TheRxFsk|Lowpass|R.ReadAddressSample\(3) & \TheRxFsk|Lowpass|R.ReadAddressSample\(2) & \TheRxFsk|Lowpass|R.ReadAddressSample[1]~DUPLICATE_q\ & \TheRxFsk|Lowpass|R.ReadAddressSample[0]~DUPLICATE_q\);

\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a0~portbdataout\ <= \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(0);
\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a1\ <= \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(1);
\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a2\ <= \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(2);
\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a3\ <= \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(3);
\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a4\ <= \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(4);
\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a5\ <= \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(5);
\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a6\ <= \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(6);
\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a7\ <= \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(7);
\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a8\ <= \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(8);
\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a9\ <= \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(9);
\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a10\ <= \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(10);
\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a11\ <= \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(11);
\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a12\ <= \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(12);
\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a13\ <= \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(13);
\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a14\ <= \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(14);
\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a15\ <= \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(15);

\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_AX_bus\ <= (\TheRxFsk|Bandpasses:7:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a15\ & \TheRxFsk|Bandpasses:7:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a15\ & 
\TheRxFsk|Bandpasses:7:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a15\ & \TheRxFsk|Bandpasses:7:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a14\ & \TheRxFsk|Bandpasses:7:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a13\ & 
\TheRxFsk|Bandpasses:7:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a12\ & \TheRxFsk|Bandpasses:7:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a11\ & \TheRxFsk|Bandpasses:7:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a10\ & 
\TheRxFsk|Bandpasses:7:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a9\ & \TheRxFsk|Bandpasses:7:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a8\ & \TheRxFsk|Bandpasses:7:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a7\ & 
\TheRxFsk|Bandpasses:7:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a6\ & \TheRxFsk|Bandpasses:7:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a5\ & \TheRxFsk|Bandpasses:7:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a4\ & 
\TheRxFsk|Bandpasses:7:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a3\ & \TheRxFsk|Bandpasses:7:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a2\ & \TheRxFsk|Bandpasses:7:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a1\ & 
\TheRxFsk|Bandpasses:7:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a0\);

\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_AY_bus\ <= (\TheRxFsk|Bandpasses:7:Bandpass1|Sample[0]~15_combout\ & \TheRxFsk|Bandpasses:7:Bandpass1|Sample[0]~15_combout\ & \TheRxFsk|Bandpasses:7:Bandpass1|Sample[0]~15_combout\ & 
\TheRxFsk|Bandpasses:7:Bandpass1|Sample[0]~15_combout\ & \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-1]~14_combout\ & \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-2]~13_combout\ & \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-3]~12_combout\ & 
\TheRxFsk|Bandpasses:7:Bandpass1|Sample[-4]~11_combout\ & \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-5]~10_combout\ & \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-6]~9_combout\ & \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-7]~8_combout\ & 
\TheRxFsk|Bandpasses:7:Bandpass1|Sample[-8]~7_combout\ & \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-9]~6_combout\ & \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-10]~5_combout\ & \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-11]~4_combout\ & 
\TheRxFsk|Bandpasses:7:Bandpass1|Sample[-12]~3_combout\ & \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-13]~2_combout\ & \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-14]~1_combout\ & \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-15]~0_combout\);

\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_resulta\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(0);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~9\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(1);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~10\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(2);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~11\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(3);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~12\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(4);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~13\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(5);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~14\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(6);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~15\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(7);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~16\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(8);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~17\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(9);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~18\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(10);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~19\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(11);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~20\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(12);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~21\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(13);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~22\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(14);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~23\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(15);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~24\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(16);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~25\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(17);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~26\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(18);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~27\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(19);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~28\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(20);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~29\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(21);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~30\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(22);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~31\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(23);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~32\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(24);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~33\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(25);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~34\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(26);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~35\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(27);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~36\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(28);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~37\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(29);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~38\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(30);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~39\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(31);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~40\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(32);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~41\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(33);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~42\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(34);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~43\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(35);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~44\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(36);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~45\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(37);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~46\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(38);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~47\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(39);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~48\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(40);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~49\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(41);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~50\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(42);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~51\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(43);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~52\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(44);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~53\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(45);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~54\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(46);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~55\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(47);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~56\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(48);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~57\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(49);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~58\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(50);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~59\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(51);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~60\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(52);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~61\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(53);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~62\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(54);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~63\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(55);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~64\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(56);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~65\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(57);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~66\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(58);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~67\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(59);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~68\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(60);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~69\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(61);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~70\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(62);
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~71\ <= \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\(63);

\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_AX_bus\ <= (\TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a15\ & \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a15\ & 
\TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a15\ & \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a14\ & \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a13\ & 
\TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a12\ & \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a11\ & \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a10\ & 
\TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a9\ & \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a8\ & \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a7\ & 
\TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a6\ & \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a5\ & \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a4~portadataout\
& \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a3\ & \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a2\ & \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a1\ & 
\TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a0~portadataout\);

\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_AY_bus\ <= (\TheRxFsk|Bandpasses:4:Bandpass1|Sample[0]~15_combout\ & \TheRxFsk|Bandpasses:4:Bandpass1|Sample[0]~15_combout\ & \TheRxFsk|Bandpasses:4:Bandpass1|Sample[0]~15_combout\ & 
\TheRxFsk|Bandpasses:4:Bandpass1|Sample[0]~15_combout\ & \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-1]~14_combout\ & \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-2]~13_combout\ & \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-3]~12_combout\ & 
\TheRxFsk|Bandpasses:4:Bandpass1|Sample[-4]~11_combout\ & \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-5]~10_combout\ & \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-6]~9_combout\ & \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-7]~8_combout\ & 
\TheRxFsk|Bandpasses:4:Bandpass1|Sample[-8]~7_combout\ & \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-9]~6_combout\ & \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-10]~5_combout\ & \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-11]~4_combout\ & 
\TheRxFsk|Bandpasses:4:Bandpass1|Sample[-12]~3_combout\ & \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-13]~2_combout\ & \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-14]~1_combout\ & \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-15]~0_combout\);

\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_resulta\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(0);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~9\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(1);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~10\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(2);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~11\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(3);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~12\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(4);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~13\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(5);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~14\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(6);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~15\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(7);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~16\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(8);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~17\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(9);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~18\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(10);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~19\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(11);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~20\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(12);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~21\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(13);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~22\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(14);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~23\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(15);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~24\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(16);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~25\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(17);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~26\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(18);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~27\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(19);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~28\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(20);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~29\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(21);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~30\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(22);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~31\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(23);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~32\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(24);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~33\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(25);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~34\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(26);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~35\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(27);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~36\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(28);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~37\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(29);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~38\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(30);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~39\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(31);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~40\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(32);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~41\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(33);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~42\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(34);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~43\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(35);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~44\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(36);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~45\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(37);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~46\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(38);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~47\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(39);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~48\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(40);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~49\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(41);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~50\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(42);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~51\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(43);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~52\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(44);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~53\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(45);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~54\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(46);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~55\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(47);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~56\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(48);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~57\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(49);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~58\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(50);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~59\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(51);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~60\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(52);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~61\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(53);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~62\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(54);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~63\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(55);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~64\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(56);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~65\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(57);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~66\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(58);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~67\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(59);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~68\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(60);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~69\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(61);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~70\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(62);
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~71\ <= \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\(63);

\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_AX_bus\ <= (\TheRxFsk|Bandpasses:7:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a15\ & \TheRxFsk|Bandpasses:7:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a15\ & 
\TheRxFsk|Bandpasses:7:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a15\ & \TheRxFsk|Bandpasses:7:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a14\ & \TheRxFsk|Bandpasses:7:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a13\ & 
\TheRxFsk|Bandpasses:7:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a12\ & \TheRxFsk|Bandpasses:7:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a11\ & \TheRxFsk|Bandpasses:7:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a10\ & 
\TheRxFsk|Bandpasses:7:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a9\ & \TheRxFsk|Bandpasses:7:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a8\ & \TheRxFsk|Bandpasses:7:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a7\ & 
\TheRxFsk|Bandpasses:7:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a6\ & \TheRxFsk|Bandpasses:7:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a5\ & \TheRxFsk|Bandpasses:7:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a4\ & 
\TheRxFsk|Bandpasses:7:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a3\ & \TheRxFsk|Bandpasses:7:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a2\ & \TheRxFsk|Bandpasses:7:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a1\ & 
\TheRxFsk|Bandpasses:7:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a0\);

\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_AY_bus\ <= (\TheRxFsk|Bandpasses:7:Bandpass0|Sample[0]~15_combout\ & \TheRxFsk|Bandpasses:7:Bandpass0|Sample[0]~15_combout\ & \TheRxFsk|Bandpasses:7:Bandpass0|Sample[0]~15_combout\ & 
\TheRxFsk|Bandpasses:7:Bandpass0|Sample[0]~15_combout\ & \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-1]~14_combout\ & \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-2]~13_combout\ & \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-3]~12_combout\ & 
\TheRxFsk|Bandpasses:7:Bandpass0|Sample[-4]~11_combout\ & \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-5]~10_combout\ & \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-6]~9_combout\ & \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-7]~8_combout\ & 
\TheRxFsk|Bandpasses:7:Bandpass0|Sample[-8]~7_combout\ & \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-9]~6_combout\ & \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-10]~5_combout\ & \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-11]~4_combout\ & 
\TheRxFsk|Bandpasses:7:Bandpass0|Sample[-12]~3_combout\ & \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-13]~2_combout\ & \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-14]~1_combout\ & \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-15]~0_combout\);

\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_resulta\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(0);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~9\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(1);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~10\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(2);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~11\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(3);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~12\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(4);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~13\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(5);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~14\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(6);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~15\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(7);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~16\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(8);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~17\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(9);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~18\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(10);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~19\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(11);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~20\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(12);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~21\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(13);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~22\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(14);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~23\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(15);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~24\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(16);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~25\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(17);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~26\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(18);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~27\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(19);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~28\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(20);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~29\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(21);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~30\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(22);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~31\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(23);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~32\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(24);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~33\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(25);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~34\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(26);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~35\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(27);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~36\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(28);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~37\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(29);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~38\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(30);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~39\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(31);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~40\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(32);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~41\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(33);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~42\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(34);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~43\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(35);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~44\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(36);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~45\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(37);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~46\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(38);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~47\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(39);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~48\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(40);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~49\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(41);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~50\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(42);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~51\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(43);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~52\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(44);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~53\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(45);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~54\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(46);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~55\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(47);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~56\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(48);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~57\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(49);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~58\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(50);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~59\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(51);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~60\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(52);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~61\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(53);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~62\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(54);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~63\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(55);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~64\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(56);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~65\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(57);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~66\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(58);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~67\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(59);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~68\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(60);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~69\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(61);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~70\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(62);
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~71\ <= \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\(63);

\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_AX_bus\ <= (\TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a15\ & \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a15\ & 
\TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a15\ & \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a14\ & \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a13\ & 
\TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a12~portadataout\ & \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a11\ & 
\TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a10\ & \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a9\ & \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a8\ & 
\TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a7\ & \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a6\ & \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a5\ & 
\TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a4\ & \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a3\ & \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a2\ & 
\TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a1\ & \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a0~portadataout\);

\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_AY_bus\ <= (\TheRxFsk|Bandpasses:4:Bandpass0|Sample[0]~15_combout\ & \TheRxFsk|Bandpasses:4:Bandpass0|Sample[0]~15_combout\ & \TheRxFsk|Bandpasses:4:Bandpass0|Sample[0]~15_combout\ & 
\TheRxFsk|Bandpasses:4:Bandpass0|Sample[0]~15_combout\ & \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-1]~14_combout\ & \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-2]~13_combout\ & \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-3]~12_combout\ & 
\TheRxFsk|Bandpasses:4:Bandpass0|Sample[-4]~11_combout\ & \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-5]~10_combout\ & \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-6]~9_combout\ & \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-7]~8_combout\ & 
\TheRxFsk|Bandpasses:4:Bandpass0|Sample[-8]~7_combout\ & \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-9]~6_combout\ & \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-10]~5_combout\ & \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-11]~4_combout\ & 
\TheRxFsk|Bandpasses:4:Bandpass0|Sample[-12]~3_combout\ & \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-13]~2_combout\ & \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-14]~1_combout\ & \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-15]~0_combout\);

\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_resulta\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(0);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~9\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(1);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~10\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(2);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~11\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(3);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~12\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(4);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~13\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(5);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~14\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(6);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~15\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(7);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~16\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(8);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~17\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(9);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~18\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(10);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~19\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(11);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~20\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(12);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~21\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(13);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~22\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(14);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~23\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(15);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~24\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(16);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~25\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(17);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~26\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(18);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~27\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(19);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~28\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(20);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~29\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(21);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~30\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(22);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~31\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(23);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~32\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(24);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~33\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(25);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~34\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(26);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~35\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(27);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~36\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(28);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~37\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(29);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~38\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(30);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~39\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(31);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~40\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(32);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~41\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(33);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~42\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(34);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~43\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(35);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~44\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(36);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~45\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(37);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~46\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(38);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~47\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(39);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~48\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(40);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~49\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(41);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~50\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(42);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~51\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(43);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~52\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(44);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~53\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(45);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~54\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(46);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~55\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(47);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~56\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(48);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~57\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(49);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~58\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(50);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~59\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(51);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~60\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(52);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~61\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(53);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~62\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(54);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~63\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(55);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~64\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(56);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~65\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(57);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~66\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(58);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~67\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(59);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~68\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(60);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~69\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(61);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~70\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(62);
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~71\ <= \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\(63);

\TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a0_PORTAADDR_bus\ <= (\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(8) & \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[7]~DUPLICATE_q\ & 
\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[6]~DUPLICATE_q\ & \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[5]~DUPLICATE_q\ & \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[4]~DUPLICATE_q\ & 
\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(3) & \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(2) & \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[1]~DUPLICATE_q\ & \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[0]~DUPLICATE_q\);

\TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a0~portadataout\ <= \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a0_PORTADATAOUT_bus\(0);
\TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a1\ <= \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a0_PORTADATAOUT_bus\(1);
\TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a2\ <= \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a0_PORTADATAOUT_bus\(2);
\TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a3\ <= \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a0_PORTADATAOUT_bus\(3);
\TheRxFsk|Bandpasses:7:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a0\ <= \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a0_PORTADATAOUT_bus\(4);
\TheRxFsk|Bandpasses:7:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a1\ <= \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a0_PORTADATAOUT_bus\(5);
\TheRxFsk|Bandpasses:7:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a2\ <= \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a0_PORTADATAOUT_bus\(6);
\TheRxFsk|Bandpasses:7:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a3\ <= \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a0_PORTADATAOUT_bus\(7);
\TheRxFsk|Bandpasses:7:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a4\ <= \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a0_PORTADATAOUT_bus\(8);
\TheRxFsk|Bandpasses:7:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a5\ <= \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a0_PORTADATAOUT_bus\(9);
\TheRxFsk|Bandpasses:7:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a6\ <= \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a0_PORTADATAOUT_bus\(10);
\TheRxFsk|Bandpasses:7:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a7\ <= \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a0_PORTADATAOUT_bus\(11);
\TheRxFsk|Bandpasses:7:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a8\ <= \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a0_PORTADATAOUT_bus\(12);
\TheRxFsk|Bandpasses:7:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a9\ <= \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a0_PORTADATAOUT_bus\(13);
\TheRxFsk|Bandpasses:7:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a10\ <= \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a0_PORTADATAOUT_bus\(14);
\TheRxFsk|Bandpasses:7:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a11\ <= \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a0_PORTADATAOUT_bus\(15);
\TheRxFsk|Bandpasses:7:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a12\ <= \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a0_PORTADATAOUT_bus\(16);
\TheRxFsk|Bandpasses:7:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a13\ <= \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a0_PORTADATAOUT_bus\(17);
\TheRxFsk|Bandpasses:7:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a14\ <= \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a0_PORTADATAOUT_bus\(18);
\TheRxFsk|Bandpasses:7:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a15\ <= \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a0_PORTADATAOUT_bus\(19);

\TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a4_PORTAADDR_bus\ <= (\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(8) & \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[7]~DUPLICATE_q\ & 
\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[6]~DUPLICATE_q\ & \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[5]~DUPLICATE_q\ & \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[4]~DUPLICATE_q\ & 
\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(3) & \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(2) & \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[1]~DUPLICATE_q\ & \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[0]~DUPLICATE_q\);

\TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a4~portadataout\ <= \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a4_PORTADATAOUT_bus\(0);
\TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a5\ <= \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a4_PORTADATAOUT_bus\(1);
\TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a6\ <= \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a4_PORTADATAOUT_bus\(2);
\TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a7\ <= \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a4_PORTADATAOUT_bus\(3);
\TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a8\ <= \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a4_PORTADATAOUT_bus\(4);
\TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a9\ <= \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a4_PORTADATAOUT_bus\(5);
\TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a10\ <= \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a4_PORTADATAOUT_bus\(6);
\TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a11\ <= \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a4_PORTADATAOUT_bus\(7);
\TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a12\ <= \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a4_PORTADATAOUT_bus\(8);
\TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a13\ <= \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a4_PORTADATAOUT_bus\(9);
\TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a14\ <= \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a4_PORTADATAOUT_bus\(10);
\TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a15\ <= \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a4_PORTADATAOUT_bus\(11);
\TheRxFsk|Bandpasses:7:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a0\ <= \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a4_PORTADATAOUT_bus\(12);
\TheRxFsk|Bandpasses:7:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a1\ <= \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a4_PORTADATAOUT_bus\(13);
\TheRxFsk|Bandpasses:7:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a2\ <= \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a4_PORTADATAOUT_bus\(14);
\TheRxFsk|Bandpasses:7:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a3\ <= \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a4_PORTADATAOUT_bus\(15);
\TheRxFsk|Bandpasses:7:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a4\ <= \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a4_PORTADATAOUT_bus\(16);
\TheRxFsk|Bandpasses:7:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a5\ <= \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a4_PORTADATAOUT_bus\(17);
\TheRxFsk|Bandpasses:7:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a6\ <= \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a4_PORTADATAOUT_bus\(18);
\TheRxFsk|Bandpasses:7:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a7\ <= \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a4_PORTADATAOUT_bus\(19);

\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTADATAIN_bus\ <= (\TheI2sToPar|D\(15) & \TheI2sToPar|D\(14) & \TheI2sToPar|D\(13) & \TheI2sToPar|D\(12) & \TheI2sToPar|D\(11) & \TheI2sToPar|D\(10) & 
\TheI2sToPar|D\(9) & \TheI2sToPar|D\(8) & \TheI2sToPar|D\(7) & \TheI2sToPar|D\(6) & \TheI2sToPar|D\(5) & \TheI2sToPar|D\(4) & \TheI2sToPar|D\(3) & \TheI2sToPar|D\(2) & \TheI2sToPar|D\(1) & \TheI2sToPar|D\(0) & \TheI2sToPar|D\(3) & 
\TheI2sToPar|D\(2) & \TheI2sToPar|D\(1) & \TheI2sToPar|D\(0));

\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTAADDR_bus\ <= (\TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[8]~_wirecell_combout\ & \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(7) & 
\TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(6) & \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[5]~DUPLICATE_q\ & \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(4) & \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(3) & 
\TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(2) & \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(1) & \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[0]~_wirecell_combout\);

\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBADDR_bus\ <= (\TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(8) & \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(7) & 
\TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(6) & \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(5) & \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(4) & \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(3) & 
\TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(2) & \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(1) & \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(0));

\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a0~portbdataout\ <= \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(0);
\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a1\ <= \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(1);
\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a2\ <= \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(2);
\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a3\ <= \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(3);
\TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a0\ <= \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(4);
\TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a1\ <= \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(5);
\TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a2\ <= \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(6);
\TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a3\ <= \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(7);
\TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a4\ <= \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(8);
\TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a5\ <= \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(9);
\TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a6\ <= \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(10);
\TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a7\ <= \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(11);
\TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a8\ <= \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(12);
\TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a9\ <= \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(13);
\TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a10\ <= \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(14);
\TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a11\ <= \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(15);
\TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a12\ <= \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(16);
\TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a13\ <= \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(17);
\TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a14\ <= \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(18);
\TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a15\ <= \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(19);

\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a4_PORTADATAIN_bus\ <= (\TheI2sToPar|D\(7) & \TheI2sToPar|D\(6) & \TheI2sToPar|D\(5) & \TheI2sToPar|D\(4) & \TheI2sToPar|D\(3) & \TheI2sToPar|D\(2) & 
\TheI2sToPar|D\(1) & \TheI2sToPar|D\(0) & \TheI2sToPar|D\(15) & \TheI2sToPar|D\(14) & \TheI2sToPar|D\(13) & \TheI2sToPar|D\(12) & \TheI2sToPar|D\(11) & \TheI2sToPar|D\(10) & \TheI2sToPar|D\(9) & \TheI2sToPar|D\(8) & \TheI2sToPar|D\(7) & 
\TheI2sToPar|D\(6) & \TheI2sToPar|D\(5) & \TheI2sToPar|D\(4));

\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a4_PORTAADDR_bus\ <= (\TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[8]~_wirecell_combout\ & \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(7) & 
\TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(6) & \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[5]~DUPLICATE_q\ & \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(4) & \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(3) & 
\TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(2) & \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(1) & \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[0]~_wirecell_combout\);

\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a4_PORTBADDR_bus\ <= (\TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(8) & \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(7) & 
\TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(6) & \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(5) & \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(4) & \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(3) & 
\TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(2) & \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(1) & \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(0));

\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a4~portbdataout\ <= \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a4_PORTBDATAOUT_bus\(0);
\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a5\ <= \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a4_PORTBDATAOUT_bus\(1);
\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a6\ <= \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a4_PORTBDATAOUT_bus\(2);
\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a7\ <= \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a4_PORTBDATAOUT_bus\(3);
\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a8\ <= \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a4_PORTBDATAOUT_bus\(4);
\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a9\ <= \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a4_PORTBDATAOUT_bus\(5);
\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a10\ <= \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a4_PORTBDATAOUT_bus\(6);
\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a11\ <= \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a4_PORTBDATAOUT_bus\(7);
\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a12\ <= \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a4_PORTBDATAOUT_bus\(8);
\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a13\ <= \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a4_PORTBDATAOUT_bus\(9);
\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a14\ <= \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a4_PORTBDATAOUT_bus\(10);
\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a15\ <= \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a4_PORTBDATAOUT_bus\(11);
\TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a0\ <= \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a4_PORTBDATAOUT_bus\(12);
\TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a1\ <= \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a4_PORTBDATAOUT_bus\(13);
\TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a2\ <= \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a4_PORTBDATAOUT_bus\(14);
\TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a3\ <= \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a4_PORTBDATAOUT_bus\(15);
\TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a4\ <= \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a4_PORTBDATAOUT_bus\(16);
\TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a5\ <= \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a4_PORTBDATAOUT_bus\(17);
\TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a6\ <= \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a4_PORTBDATAOUT_bus\(18);
\TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a7\ <= \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a4_PORTBDATAOUT_bus\(19);

\TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a0_PORTAADDR_bus\ <= (\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(8) & \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[7]~DUPLICATE_q\ & 
\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[6]~DUPLICATE_q\ & \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[5]~DUPLICATE_q\ & \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[4]~DUPLICATE_q\ & 
\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(3) & \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(2) & \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[1]~DUPLICATE_q\ & \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[0]~DUPLICATE_q\);

\TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a0~portadataout\ <= \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a0_PORTADATAOUT_bus\(0);
\TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a1\ <= \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a0_PORTADATAOUT_bus\(1);
\TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a2\ <= \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a0_PORTADATAOUT_bus\(2);
\TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a3\ <= \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a0_PORTADATAOUT_bus\(3);
\TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a4\ <= \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a0_PORTADATAOUT_bus\(4);
\TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a5\ <= \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a0_PORTADATAOUT_bus\(5);
\TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a6\ <= \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a0_PORTADATAOUT_bus\(6);
\TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a7\ <= \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a0_PORTADATAOUT_bus\(7);
\TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a8\ <= \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a0_PORTADATAOUT_bus\(8);
\TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a9\ <= \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a0_PORTADATAOUT_bus\(9);
\TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a10\ <= \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a0_PORTADATAOUT_bus\(10);
\TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a11\ <= \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a0_PORTADATAOUT_bus\(11);
\TheRxFsk|Bandpasses:7:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a8\ <= \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a0_PORTADATAOUT_bus\(12);
\TheRxFsk|Bandpasses:7:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a9\ <= \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a0_PORTADATAOUT_bus\(13);
\TheRxFsk|Bandpasses:7:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a10\ <= \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a0_PORTADATAOUT_bus\(14);
\TheRxFsk|Bandpasses:7:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a11\ <= \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a0_PORTADATAOUT_bus\(15);
\TheRxFsk|Bandpasses:7:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a12\ <= \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a0_PORTADATAOUT_bus\(16);
\TheRxFsk|Bandpasses:7:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a13\ <= \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a0_PORTADATAOUT_bus\(17);
\TheRxFsk|Bandpasses:7:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a14\ <= \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a0_PORTADATAOUT_bus\(18);
\TheRxFsk|Bandpasses:7:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a15\ <= \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a0_PORTADATAOUT_bus\(19);

\TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a12_PORTAADDR_bus\ <= (\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(8) & \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[7]~DUPLICATE_q\ & 
\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[6]~DUPLICATE_q\ & \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[5]~DUPLICATE_q\ & \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[4]~DUPLICATE_q\ & 
\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(3) & \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(2) & \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[1]~DUPLICATE_q\ & \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[0]~DUPLICATE_q\);

\TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a12~portadataout\ <= \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a12_PORTADATAOUT_bus\(0);
\TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a13\ <= \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a12_PORTADATAOUT_bus\(1);
\TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a14\ <= \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a12_PORTADATAOUT_bus\(2);
\TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a15\ <= \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a12_PORTADATAOUT_bus\(3);

\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTADATAIN_bus\ <= (\TheI2sToPar|D\(15) & \TheI2sToPar|D\(14) & \TheI2sToPar|D\(13) & \TheI2sToPar|D\(12) & \TheI2sToPar|D\(11) & \TheI2sToPar|D\(10) & 
\TheI2sToPar|D\(9) & \TheI2sToPar|D\(8) & \TheI2sToPar|D\(11) & \TheI2sToPar|D\(10) & \TheI2sToPar|D\(9) & \TheI2sToPar|D\(8) & \TheI2sToPar|D\(7) & \TheI2sToPar|D\(6) & \TheI2sToPar|D\(5) & \TheI2sToPar|D\(4) & \TheI2sToPar|D\(3) & 
\TheI2sToPar|D\(2) & \TheI2sToPar|D\(1) & \TheI2sToPar|D\(0));

\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTAADDR_bus\ <= (\TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[8]~_wirecell_combout\ & \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(7) & 
\TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(6) & \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[5]~DUPLICATE_q\ & \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(4) & \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(3) & 
\TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(2) & \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(1) & \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[0]~_wirecell_combout\);

\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBADDR_bus\ <= (\TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(8) & \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(7) & 
\TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(6) & \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(5) & \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(4) & \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(3) & 
\TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(2) & \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(1) & \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(0));

\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a0~portbdataout\ <= \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(0);
\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a1\ <= \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(1);
\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a2\ <= \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(2);
\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a3\ <= \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(3);
\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a4\ <= \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(4);
\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a5\ <= \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(5);
\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a6\ <= \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(6);
\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a7\ <= \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(7);
\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a8\ <= \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(8);
\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a9\ <= \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(9);
\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a10\ <= \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(10);
\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a11\ <= \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(11);
\TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a8\ <= \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(12);
\TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a9\ <= \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(13);
\TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a10\ <= \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(14);
\TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a11\ <= \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(15);
\TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a12\ <= \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(16);
\TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a13\ <= \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(17);
\TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a14\ <= \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(18);
\TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a15\ <= \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\(19);

\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a12_PORTADATAIN_bus\ <= (gnd & gnd & gnd & gnd & gnd & gnd & gnd & gnd & gnd & gnd & gnd & gnd & gnd & gnd & gnd & gnd & \TheI2sToPar|D\(15) & \TheI2sToPar|D\(14) & 
\TheI2sToPar|D\(13) & \TheI2sToPar|D\(12));

\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a12_PORTAADDR_bus\ <= (\TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[8]~_wirecell_combout\ & \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(7) & 
\TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(6) & \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[5]~DUPLICATE_q\ & \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(4) & \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(3) & 
\TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(2) & \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(1) & \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[0]~_wirecell_combout\);

\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a12_PORTBADDR_bus\ <= (\TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(8) & \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(7) & 
\TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(6) & \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(5) & \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(4) & \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(3) & 
\TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(2) & \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(1) & \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(0));

\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a12~portbdataout\ <= \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a12_PORTBDATAOUT_bus\(0);
\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a13\ <= \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a12_PORTBDATAOUT_bus\(1);
\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a14\ <= \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a12_PORTBDATAOUT_bus\(2);
\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a15\ <= \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a12_PORTBDATAOUT_bus\(3);

\PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_VCOPH0\ <= \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_VCOPH_bus\(0);
\PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_VCOPH1\ <= \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_VCOPH_bus\(1);
\PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_VCOPH2\ <= \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_VCOPH_bus\(2);
\PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_VCOPH3\ <= \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_VCOPH_bus\(3);
\PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_VCOPH4\ <= \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_VCOPH_bus\(4);
\PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_VCOPH5\ <= \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_VCOPH_bus\(5);
\PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_VCOPH6\ <= \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_VCOPH_bus\(6);
\PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_VCOPH7\ <= \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_VCOPH_bus\(7);

\PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_MHI0\ <= \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_MHI_bus\(0);
\PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_MHI1\ <= \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_MHI_bus\(1);
\PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_MHI2\ <= \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_MHI_bus\(2);
\PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_MHI3\ <= \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_MHI_bus\(3);
\PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_MHI4\ <= \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_MHI_bus\(4);
\PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_MHI5\ <= \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_MHI_bus\(5);
\PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_MHI6\ <= \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_MHI_bus\(6);
\PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_MHI7\ <= \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_MHI_bus\(7);

\PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~PLL_REFCLK_SELECT_CLKIN_bus\ <= (gnd & gnd & gnd & \iClk~input_o\);

\PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~PLL_RECONFIG_MHI_bus\ <= (
\PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_MHI7\ & 
\PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_MHI6\ & 
\PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_MHI5\ & 
\PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_MHI4\ & 
\PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_MHI3\ & 
\PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_MHI2\ & 
\PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_MHI1\ & 
\PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_MHI0\);

\PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~PLL_RECONFIGSHIFTEN6\ <= \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~PLL_RECONFIG_SHIFTEN_bus\(6);

\PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~PLL_OUTPUT_COUNTER_VCO0PH_bus\ <= (
\PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_VCOPH7\ & 
\PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_VCOPH6\ & 
\PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_VCOPH5\ & 
\PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_VCOPH4\ & 
\PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_VCOPH3\ & 
\PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_VCOPH2\ & 
\PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_VCOPH1\ & 
\PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_VCOPH0\);
\TheRxFsk|ALT_INV_Add2~37_sumout\ <= NOT \TheRxFsk|Add2~37_sumout\;
\TheRxFsk|ALT_INV_Add2~33_sumout\ <= NOT \TheRxFsk|Add2~33_sumout\;
\TheRxFsk|ALT_INV_Add2~29_sumout\ <= NOT \TheRxFsk|Add2~29_sumout\;
\TheRxFsk|ALT_INV_Add2~25_sumout\ <= NOT \TheRxFsk|Add2~25_sumout\;
\TheRxFsk|ALT_INV_Add2~21_sumout\ <= NOT \TheRxFsk|Add2~21_sumout\;
\TheRxFsk|ALT_INV_Add2~17_sumout\ <= NOT \TheRxFsk|Add2~17_sumout\;
\TheRxFsk|ALT_INV_Add2~13_sumout\ <= NOT \TheRxFsk|Add2~13_sumout\;
\TheRxFsk|ALT_INV_Add2~9_sumout\ <= NOT \TheRxFsk|Add2~9_sumout\;
\TheRxFsk|ALT_INV_Add2~5_sumout\ <= NOT \TheRxFsk|Add2~5_sumout\;
\TheRxFsk|ALT_INV_Add2~1_sumout\ <= NOT \TheRxFsk|Add2~1_sumout\;
\TheRxFsk|Lowpass|ALT_INV_Add4~17_sumout\ <= NOT \TheRxFsk|Lowpass|Add4~17_sumout\;
\TheRxFsk|Lowpass|ALT_INV_Sum[-2]~q\ <= NOT \TheRxFsk|Lowpass|Sum[-2]~q\;
\TheRxFsk|Lowpass|ALT_INV_DdryDelayed\(0) <= NOT \TheRxFsk|Lowpass|DdryDelayed\(0);
\TheRxFsk|Lowpass|ALT_INV_DdryDelayed[-1]~q\ <= NOT \TheRxFsk|Lowpass|DdryDelayed[-1]~q\;
\TheRxFsk|Lowpass|ALT_INV_DdryDelayed[-2]~q\ <= NOT \TheRxFsk|Lowpass|DdryDelayed[-2]~q\;
\TheRxFsk|Lowpass|ALT_INV_DdryDelayed[-3]~q\ <= NOT \TheRxFsk|Lowpass|DdryDelayed[-3]~q\;
\TheRxFsk|Lowpass|ALT_INV_DdryDelayed[-4]~q\ <= NOT \TheRxFsk|Lowpass|DdryDelayed[-4]~q\;
\TheRxFsk|Lowpass|ALT_INV_DdryDelayed[-5]~q\ <= NOT \TheRxFsk|Lowpass|DdryDelayed[-5]~q\;
\TheRxFsk|Lowpass|ALT_INV_DdryDelayed[-6]~q\ <= NOT \TheRxFsk|Lowpass|DdryDelayed[-6]~q\;
\TheRxFsk|Lowpass|ALT_INV_DdryDelayed[-7]~q\ <= NOT \TheRxFsk|Lowpass|DdryDelayed[-7]~q\;
\TheRxFsk|Lowpass|ALT_INV_DdryDelayed[-8]~q\ <= NOT \TheRxFsk|Lowpass|DdryDelayed[-8]~q\;
\TheRxFsk|Lowpass|ALT_INV_DdryDelayed[-9]~q\ <= NOT \TheRxFsk|Lowpass|DdryDelayed[-9]~q\;
\TheRxFsk|Lowpass|ALT_INV_DdryDelayed[-10]~q\ <= NOT \TheRxFsk|Lowpass|DdryDelayed[-10]~q\;
\TheRxFsk|Lowpass|ALT_INV_DdryDelayed[-11]~q\ <= NOT \TheRxFsk|Lowpass|DdryDelayed[-11]~q\;
\TheRxFsk|Lowpass|ALT_INV_DdryDelayed[-12]~q\ <= NOT \TheRxFsk|Lowpass|DdryDelayed[-12]~q\;
\TheRxFsk|Lowpass|ALT_INV_DdryDelayed[-13]~q\ <= NOT \TheRxFsk|Lowpass|DdryDelayed[-13]~q\;
\TheRxFsk|Lowpass|ALT_INV_DdryDelayed[-14]~q\ <= NOT \TheRxFsk|Lowpass|DdryDelayed[-14]~q\;
\TheRxFsk|Lowpass|ALT_INV_DdryDelayed[-15]~q\ <= NOT \TheRxFsk|Lowpass|DdryDelayed[-15]~q\;
\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a1\ <= NOT \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a1\;
\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a2\ <= NOT \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a2\;
\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a3\ <= NOT \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a3\;
\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a4\ <= NOT \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a4\;
\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a5\ <= NOT \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a5\;
\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a6\ <= NOT \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a6\;
\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a7\ <= NOT \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a7\;
\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a8\ <= NOT \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a8\;
\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a9\ <= NOT \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a9\;
\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a10\ <= NOT \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a10\;
\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a11\ <= NOT \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a11\;
\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a12\ <= NOT \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a12\;
\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a13\ <= NOT \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a13\;
\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a14\ <= NOT \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a14\;
\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a15\ <= NOT \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a15\;
\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a0~portbdataout\ <= NOT \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a0~portbdataout\;
\TheRxFsk|Lowpass|ALT_INV_Add4~13_sumout\ <= NOT \TheRxFsk|Lowpass|Add4~13_sumout\;
\TheRxFsk|Lowpass|ALT_INV_Sum[-1]~q\ <= NOT \TheRxFsk|Lowpass|Sum[-1]~q\;
\TheRxFsk|Lowpass|ALT_INV_Mult0~39\ <= NOT \TheRxFsk|Lowpass|Mult0~39\;
\TheRxFsk|Lowpass|ALT_INV_Mult0~38\ <= NOT \TheRxFsk|Lowpass|Mult0~38\;
\TheRxFsk|Lowpass|ALT_INV_Mult0~37\ <= NOT \TheRxFsk|Lowpass|Mult0~37\;
\TheRxFsk|Lowpass|ALT_INV_Mult0~36\ <= NOT \TheRxFsk|Lowpass|Mult0~36\;
\TheRxFsk|Lowpass|ALT_INV_Mult0~35\ <= NOT \TheRxFsk|Lowpass|Mult0~35\;
\TheRxFsk|Lowpass|ALT_INV_Mult0~34\ <= NOT \TheRxFsk|Lowpass|Mult0~34\;
\TheRxFsk|Lowpass|ALT_INV_Mult0~33\ <= NOT \TheRxFsk|Lowpass|Mult0~33\;
\TheRxFsk|Lowpass|ALT_INV_Mult0~32\ <= NOT \TheRxFsk|Lowpass|Mult0~32\;
\TheRxFsk|Lowpass|ALT_INV_Mult0~31\ <= NOT \TheRxFsk|Lowpass|Mult0~31\;
\TheRxFsk|Lowpass|ALT_INV_Mult0~30\ <= NOT \TheRxFsk|Lowpass|Mult0~30\;
\TheRxFsk|Lowpass|ALT_INV_Mult0~29\ <= NOT \TheRxFsk|Lowpass|Mult0~29\;
\TheRxFsk|Lowpass|ALT_INV_Mult0~28\ <= NOT \TheRxFsk|Lowpass|Mult0~28\;
\TheRxFsk|Lowpass|ALT_INV_Mult0~27\ <= NOT \TheRxFsk|Lowpass|Mult0~27\;
\TheRxFsk|Lowpass|ALT_INV_Mult0~26\ <= NOT \TheRxFsk|Lowpass|Mult0~26\;
\TheRxFsk|Lowpass|ALT_INV_Mult0~25\ <= NOT \TheRxFsk|Lowpass|Mult0~25\;
\TheRxFsk|Lowpass|ALT_INV_Mult0~24\ <= NOT \TheRxFsk|Lowpass|Mult0~24\;
\TheRxFsk|Lowpass|ALT_INV_Mult0~23\ <= NOT \TheRxFsk|Lowpass|Mult0~23\;
\TheRxFsk|Lowpass|ALT_INV_Mult0~22\ <= NOT \TheRxFsk|Lowpass|Mult0~22\;
\TheRxFsk|Lowpass|ALT_INV_Mult0~21\ <= NOT \TheRxFsk|Lowpass|Mult0~21\;
\TheRxFsk|Lowpass|ALT_INV_Mult0~20\ <= NOT \TheRxFsk|Lowpass|Mult0~20\;
\TheRxFsk|Lowpass|ALT_INV_Mult0~19\ <= NOT \TheRxFsk|Lowpass|Mult0~19\;
\TheRxFsk|Lowpass|ALT_INV_Mult0~18\ <= NOT \TheRxFsk|Lowpass|Mult0~18\;
\TheRxFsk|Lowpass|ALT_INV_Mult0~17\ <= NOT \TheRxFsk|Lowpass|Mult0~17\;
\TheRxFsk|Lowpass|ALT_INV_Mult0~16\ <= NOT \TheRxFsk|Lowpass|Mult0~16\;
\TheRxFsk|Lowpass|ALT_INV_Mult0~15\ <= NOT \TheRxFsk|Lowpass|Mult0~15\;
\TheRxFsk|Lowpass|ALT_INV_Mult0~14\ <= NOT \TheRxFsk|Lowpass|Mult0~14\;
\TheRxFsk|Lowpass|ALT_INV_Mult0~13\ <= NOT \TheRxFsk|Lowpass|Mult0~13\;
\TheRxFsk|Lowpass|ALT_INV_Mult0~12\ <= NOT \TheRxFsk|Lowpass|Mult0~12\;
\TheRxFsk|Lowpass|ALT_INV_Mult0~11\ <= NOT \TheRxFsk|Lowpass|Mult0~11\;
\TheRxFsk|Lowpass|ALT_INV_Mult0~10\ <= NOT \TheRxFsk|Lowpass|Mult0~10\;
\TheRxFsk|Lowpass|ALT_INV_Mult0~9\ <= NOT \TheRxFsk|Lowpass|Mult0~9\;
\TheRxFsk|Lowpass|ALT_INV_Mult0~8_resulta\ <= NOT \TheRxFsk|Lowpass|Mult0~8_resulta\;
\TheRxFsk|Lowpass|ALT_INV_Add2~25_sumout\ <= NOT \TheRxFsk|Lowpass|Add2~25_sumout\;
\TheRxFsk|Lowpass|ALT_INV_Add2~21_sumout\ <= NOT \TheRxFsk|Lowpass|Add2~21_sumout\;
\TheRxFsk|Lowpass|ALT_INV_Add2~13_sumout\ <= NOT \TheRxFsk|Lowpass|Add2~13_sumout\;
\TheRxFsk|Lowpass|ALT_INV_Add2~9_sumout\ <= NOT \TheRxFsk|Lowpass|Add2~9_sumout\;
\TheRxFsk|Lowpass|ALT_INV_Add2~5_sumout\ <= NOT \TheRxFsk|Lowpass|Add2~5_sumout\;
\TheRxFsk|Lowpass|ALT_INV_Add2~1_sumout\ <= NOT \TheRxFsk|Lowpass|Add2~1_sumout\;
\TheRxFsk|Lowpass|ALT_INV_Add4~9_sumout\ <= NOT \TheRxFsk|Lowpass|Add4~9_sumout\;
\TheRxFsk|Lowpass|ALT_INV_Add3~1_sumout\ <= NOT \TheRxFsk|Lowpass|Add3~1_sumout\;
\TheRxFsk|Lowpass|ALT_INV_Add4~5_sumout\ <= NOT \TheRxFsk|Lowpass|Add4~5_sumout\;
\GenClks|ALT_INV_Add0~29_sumout\ <= NOT \GenClks|Add0~29_sumout\;
\GenClks|ALT_INV_Add0~13_sumout\ <= NOT \GenClks|Add0~13_sumout\;
\TheRxFsk|Lowpass|ALT_INV_Add4~1_sumout\ <= NOT \TheRxFsk|Lowpass|Add4~1_sumout\;
\TheRxFsk|Lowpass|ALT_INV_Sum\(0) <= NOT \TheRxFsk|Lowpass|Sum\(0);
\ConfigureCodec|ALT_INV_R.AddrCtr\(0) <= NOT \ConfigureCodec|R.AddrCtr\(0);
\ConfigureCodec|ALT_INV_R.AddrCtr\(3) <= NOT \ConfigureCodec|R.AddrCtr\(3);
\ConfigureCodec|ALT_INV_R.AddrCtr\(4) <= NOT \ConfigureCodec|R.AddrCtr\(4);
\ConfigureCodec|ALT_INV_R.AddrCtr\(5) <= NOT \ConfigureCodec|R.AddrCtr\(5);
\ConfigureCodec|ALT_INV_R.AddrCtr\(6) <= NOT \ConfigureCodec|R.AddrCtr\(6);
\ConfigureCodec|ALT_INV_R.AddrCtr\(1) <= NOT \ConfigureCodec|R.AddrCtr\(1);
\ConfigureCodec|ALT_INV_R.AddrCtr\(2) <= NOT \ConfigureCodec|R.AddrCtr\(2);
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.EnableSumUp~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|R.EnableSumUp~q\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.SelSumUp~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|R.SelSumUp~q\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_R.EnableSumUp~q\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|R.EnableSumUp~q\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_R.SelSumUp~q\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|R.SelSumUp~q\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_R.EnableSumUp~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|R.EnableSumUp~q\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_R.SelSumUp~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|R.SelSumUp~q\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_R.EnableSumUp~q\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|R.EnableSumUp~q\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_R.SelSumUp~q\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|R.SelSumUp~q\;
\TheRxFsk|Lowpass|ALT_INV_MultResult[-4]~3_combout\ <= NOT \TheRxFsk|Lowpass|MultResult[-4]~3_combout\;
\TheRxFsk|ALT_INV_Mux1~0_combout\ <= NOT \TheRxFsk|Mux1~0_combout\;
\TheRxFsk|ALT_INV_Mux17~0_combout\ <= NOT \TheRxFsk|Mux17~0_combout\;
\TheRxFsk|ALT_INV_Mux2~0_combout\ <= NOT \TheRxFsk|Mux2~0_combout\;
\TheRxFsk|ALT_INV_Mux18~0_combout\ <= NOT \TheRxFsk|Mux18~0_combout\;
\TheRxFsk|ALT_INV_Mux3~0_combout\ <= NOT \TheRxFsk|Mux3~0_combout\;
\TheRxFsk|ALT_INV_Mux19~0_combout\ <= NOT \TheRxFsk|Mux19~0_combout\;
\TheRxFsk|ALT_INV_Mux4~0_combout\ <= NOT \TheRxFsk|Mux4~0_combout\;
\TheRxFsk|ALT_INV_Mux20~0_combout\ <= NOT \TheRxFsk|Mux20~0_combout\;
\TheRxFsk|ALT_INV_Mux5~0_combout\ <= NOT \TheRxFsk|Mux5~0_combout\;
\TheRxFsk|ALT_INV_Mux21~0_combout\ <= NOT \TheRxFsk|Mux21~0_combout\;
\TheRxFsk|ALT_INV_Mux6~0_combout\ <= NOT \TheRxFsk|Mux6~0_combout\;
\TheRxFsk|ALT_INV_Mux22~0_combout\ <= NOT \TheRxFsk|Mux22~0_combout\;
\TheRxFsk|ALT_INV_Mux7~0_combout\ <= NOT \TheRxFsk|Mux7~0_combout\;
\TheRxFsk|ALT_INV_Mux23~0_combout\ <= NOT \TheRxFsk|Mux23~0_combout\;
\TheRxFsk|ALT_INV_Mux8~0_combout\ <= NOT \TheRxFsk|Mux8~0_combout\;
\TheRxFsk|ALT_INV_Mux24~0_combout\ <= NOT \TheRxFsk|Mux24~0_combout\;
\TheRxFsk|ALT_INV_Mux9~0_combout\ <= NOT \TheRxFsk|Mux9~0_combout\;
\TheRxFsk|ALT_INV_Mux25~0_combout\ <= NOT \TheRxFsk|Mux25~0_combout\;
\TheRxFsk|ALT_INV_Mux10~0_combout\ <= NOT \TheRxFsk|Mux10~0_combout\;
\TheRxFsk|ALT_INV_Mux26~0_combout\ <= NOT \TheRxFsk|Mux26~0_combout\;
\TheRxFsk|ALT_INV_Mux11~0_combout\ <= NOT \TheRxFsk|Mux11~0_combout\;
\TheRxFsk|ALT_INV_Mux27~0_combout\ <= NOT \TheRxFsk|Mux27~0_combout\;
\TheRxFsk|ALT_INV_Mux12~0_combout\ <= NOT \TheRxFsk|Mux12~0_combout\;
\TheRxFsk|ALT_INV_Mux28~0_combout\ <= NOT \TheRxFsk|Mux28~0_combout\;
\TheRxFsk|ALT_INV_Mux13~0_combout\ <= NOT \TheRxFsk|Mux13~0_combout\;
\TheRxFsk|ALT_INV_Mux29~0_combout\ <= NOT \TheRxFsk|Mux29~0_combout\;
\TheRxFsk|ALT_INV_Mux14~0_combout\ <= NOT \TheRxFsk|Mux14~0_combout\;
\TheRxFsk|ALT_INV_Mux30~0_combout\ <= NOT \TheRxFsk|Mux30~0_combout\;
\TheRxFsk|ALT_INV_Mux15~0_combout\ <= NOT \TheRxFsk|Mux15~0_combout\;
\TheRxFsk|ALT_INV_Mux31~0_combout\ <= NOT \TheRxFsk|Mux31~0_combout\;
\TheRxFsk|Bandpasses:11:Bandpass0|ALT_INV_R.SumState.Idle~q\ <= NOT \TheRxFsk|Bandpasses:11:Bandpass0|R.SumState.Idle~q\;
\TheRxFsk|Lowpass|ALT_INV_MultResult[-3]~2_combout\ <= NOT \TheRxFsk|Lowpass|MultResult[-3]~2_combout\;
\TheRxFsk|Lowpass|ALT_INV_Equal0~0_combout\ <= NOT \TheRxFsk|Lowpass|Equal0~0_combout\;
\TheRxFsk|Lowpass|ALT_INV_Equal2~0_combout\ <= NOT \TheRxFsk|Lowpass|Equal2~0_combout\;
\TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.AddressState~q\ <= NOT \TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~q\;
\TheRxFsk|Bandpasses:11:Bandpass0|ALT_INV_R.SumState.SumEnable~q\ <= NOT \TheRxFsk|Bandpasses:11:Bandpass0|R.SumState.SumEnable~q\;
\TheRxFsk|Lowpass|ALT_INV_MultResult[-2]~1_combout\ <= NOT \TheRxFsk|Lowpass|MultResult[-2]~1_combout\;
\TheRxFsk|Lowpass|ALT_INV_R.ReadAddressSample\(6) <= NOT \TheRxFsk|Lowpass|R.ReadAddressSample\(6);
\TheRxFsk|Lowpass|ALT_INV_R.ReadAddressSample\(5) <= NOT \TheRxFsk|Lowpass|R.ReadAddressSample\(5);
\TheRxFsk|Lowpass|ALT_INV_R.ReadAddressSample\(4) <= NOT \TheRxFsk|Lowpass|R.ReadAddressSample\(4);
\TheRxFsk|Lowpass|ALT_INV_R.ReadAddressSample\(3) <= NOT \TheRxFsk|Lowpass|R.ReadAddressSample\(3);
\TheRxFsk|Lowpass|ALT_INV_R.ReadAddressSample\(2) <= NOT \TheRxFsk|Lowpass|R.ReadAddressSample\(2);
\TheRxFsk|Lowpass|ALT_INV_R.ReadAddressSample\(1) <= NOT \TheRxFsk|Lowpass|R.ReadAddressSample\(1);
\TheRxFsk|Lowpass|ALT_INV_R.ReadAddressSample\(0) <= NOT \TheRxFsk|Lowpass|R.ReadAddressSample\(0);
\TheRxFsk|Lowpass|ALT_INV_R.WriteAddress\(6) <= NOT \TheRxFsk|Lowpass|R.WriteAddress\(6);
\TheRxFsk|Lowpass|ALT_INV_R.WriteAddress\(5) <= NOT \TheRxFsk|Lowpass|R.WriteAddress\(5);
\TheRxFsk|Lowpass|ALT_INV_R.WriteAddress\(4) <= NOT \TheRxFsk|Lowpass|R.WriteAddress\(4);
\TheRxFsk|Lowpass|ALT_INV_R.WriteAddress\(3) <= NOT \TheRxFsk|Lowpass|R.WriteAddress\(3);
\TheRxFsk|Lowpass|ALT_INV_R.WriteAddress\(2) <= NOT \TheRxFsk|Lowpass|R.WriteAddress\(2);
\TheRxFsk|Lowpass|ALT_INV_R.WriteAddress\(1) <= NOT \TheRxFsk|Lowpass|R.WriteAddress\(1);
\TheRxFsk|Lowpass|ALT_INV_R.WriteAddress\(0) <= NOT \TheRxFsk|Lowpass|R.WriteAddress\(0);
\TheRxFsk|Lowpass|ALT_INV_CoefMemory~7_combout\ <= NOT \TheRxFsk|Lowpass|CoefMemory~7_combout\;
\TheRxFsk|Lowpass|ALT_INV_CoefMemory~5_combout\ <= NOT \TheRxFsk|Lowpass|CoefMemory~5_combout\;
\TheRxFsk|Lowpass|ALT_INV_CoefMemory~4_combout\ <= NOT \TheRxFsk|Lowpass|CoefMemory~4_combout\;
\TheRxFsk|Lowpass|ALT_INV_CoefMemory~2_combout\ <= NOT \TheRxFsk|Lowpass|CoefMemory~2_combout\;
\TheRxFsk|Lowpass|ALT_INV_CoefMemory~1_combout\ <= NOT \TheRxFsk|Lowpass|CoefMemory~1_combout\;
\TheRxFsk|Bandpasses:11:Bandpass1|ALT_INV_Equal1~1_combout\ <= NOT \TheRxFsk|Bandpasses:11:Bandpass1|Equal1~1_combout\;
\TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.ReadAddressCoef\(0) <= NOT \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(0);
\TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.ReadAddressCoef\(1) <= NOT \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(1);
\TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.ReadAddressCoef\(2) <= NOT \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(2);
\TheRxFsk|Bandpasses:11:Bandpass1|ALT_INV_Equal1~0_combout\ <= NOT \TheRxFsk|Bandpasses:11:Bandpass1|Equal1~0_combout\;
\TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.ReadAddressCoef\(3) <= NOT \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(3);
\TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.ReadAddressCoef\(4) <= NOT \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(4);
\TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.ReadAddressCoef\(5) <= NOT \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(5);
\TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.ReadAddressCoef\(6) <= NOT \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(6);
\TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.ReadAddressCoef\(7) <= NOT \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(7);
\TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.ReadAddressCoef\(8) <= NOT \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(8);
\TheRxFsk|Bandpasses:11:Bandpass0|ALT_INV_R.SumState.SumSelect~q\ <= NOT \TheRxFsk|Bandpasses:11:Bandpass0|R.SumState.SumSelect~q\;
\TheRxFsk|Lowpass|ALT_INV_MultResult[-1]~0_combout\ <= NOT \TheRxFsk|Lowpass|MultResult[-1]~0_combout\;
\TheRxFsk|Lowpass|ALT_INV_R.FirstSample~q\ <= NOT \TheRxFsk|Lowpass|R.FirstSample~q\;
\TheRxFsk|Lowpass|ALT_INV_R.AddressState~q\ <= NOT \TheRxFsk|Lowpass|R.AddressState~q\;
\TheRxFsk|Bandpasses:11:Bandpass0|ALT_INV_R.SumState.SumWait2~q\ <= NOT \TheRxFsk|Bandpasses:11:Bandpass0|R.SumState.SumWait2~q\;
\TheRxFsk|Bandpasses:11:Bandpass0|ALT_INV_R.SumState.SumValid~q\ <= NOT \TheRxFsk|Bandpasses:11:Bandpass0|R.SumState.SumValid~q\;
\TheRxFsk|Lowpass|ALT_INV_Equal1~0_combout\ <= NOT \TheRxFsk|Lowpass|Equal1~0_combout\;
\TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(2) <= NOT \TheRxFsk|Lowpass|R.ReadAddressCoef\(2);
\TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(3) <= NOT \TheRxFsk|Lowpass|R.ReadAddressCoef\(3);
\TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(0) <= NOT \TheRxFsk|Lowpass|R.ReadAddressCoef\(0);
\TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(1) <= NOT \TheRxFsk|Lowpass|R.ReadAddressCoef\(1);
\TheRxFsk|Lowpass|ALT_INV_R.SumState.SumSelect~q\ <= NOT \TheRxFsk|Lowpass|R.SumState.SumSelect~q\;
\TheRxFsk|Lowpass|ALT_INV_CoefMemory~0_combout\ <= NOT \TheRxFsk|Lowpass|CoefMemory~0_combout\;
\TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(4) <= NOT \TheRxFsk|Lowpass|R.ReadAddressCoef\(4);
\TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(5) <= NOT \TheRxFsk|Lowpass|R.ReadAddressCoef\(5);
\TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(6) <= NOT \TheRxFsk|Lowpass|R.ReadAddressCoef\(6);
\ConfigureCodec|ALT_INV_Selector13~2_combout\ <= NOT \ConfigureCodec|Selector13~2_combout\;
\ConfigureCodec|ALT_INV_Selector12~1_combout\ <= NOT \ConfigureCodec|Selector12~1_combout\;
\ConfigureCodec|ALT_INV_Selector12~0_combout\ <= NOT \ConfigureCodec|Selector12~0_combout\;
\ConfigureCodec|ALT_INV_Selector11~2_combout\ <= NOT \ConfigureCodec|Selector11~2_combout\;
\ConfigureCodec|ALT_INV_NextR~10_combout\ <= NOT \ConfigureCodec|NextR~10_combout\;
\ConfigureCodec|ALT_INV_Mux8~0_combout\ <= NOT \ConfigureCodec|Mux8~0_combout\;
\ConfigureCodec|ALT_INV_Selector11~1_combout\ <= NOT \ConfigureCodec|Selector11~1_combout\;
\ConfigureCodec|ALT_INV_Selector11~0_combout\ <= NOT \ConfigureCodec|Selector11~0_combout\;
\ConfigureCodec|ALT_INV_Selector10~1_combout\ <= NOT \ConfigureCodec|Selector10~1_combout\;
\ConfigureCodec|ALT_INV_Selector5~0_combout\ <= NOT \ConfigureCodec|Selector5~0_combout\;
\ConfigureCodec|ALT_INV_Selector10~0_combout\ <= NOT \ConfigureCodec|Selector10~0_combout\;
\ConfigureCodec|ALT_INV_Selector13~1_combout\ <= NOT \ConfigureCodec|Selector13~1_combout\;
\ConfigureCodec|ALT_INV_Selector1~0_combout\ <= NOT \ConfigureCodec|Selector1~0_combout\;
\ConfigureCodec|ALT_INV_Selector15~2_combout\ <= NOT \ConfigureCodec|Selector15~2_combout\;
\ConfigureCodec|ALT_INV_Selector15~1_combout\ <= NOT \ConfigureCodec|Selector15~1_combout\;
\ConfigureCodec|ALT_INV_R.FrameState.Start~q\ <= NOT \ConfigureCodec|R.FrameState.Start~q\;
\ConfigureCodec|ALT_INV_Selector15~0_combout\ <= NOT \ConfigureCodec|Selector15~0_combout\;
\ConfigureCodec|ALT_INV_R.FrameState.Address~q\ <= NOT \ConfigureCodec|R.FrameState.Address~q\;
\ConfigureCodec|ALT_INV_Mux9~4_combout\ <= NOT \ConfigureCodec|Mux9~4_combout\;
\ConfigureCodec|ALT_INV_Mux9~3_combout\ <= NOT \ConfigureCodec|Mux9~3_combout\;
\ConfigureCodec|ALT_INV_R.Data\(15) <= NOT \ConfigureCodec|R.Data\(15);
\ConfigureCodec|ALT_INV_R.Data\(7) <= NOT \ConfigureCodec|R.Data\(7);
\ConfigureCodec|ALT_INV_R.Data\(11) <= NOT \ConfigureCodec|R.Data\(11);
\ConfigureCodec|ALT_INV_R.Data\(3) <= NOT \ConfigureCodec|R.Data\(3);
\ConfigureCodec|ALT_INV_Mux9~2_combout\ <= NOT \ConfigureCodec|Mux9~2_combout\;
\ConfigureCodec|ALT_INV_R.Data\(13) <= NOT \ConfigureCodec|R.Data\(13);
\ConfigureCodec|ALT_INV_R.Data\(5) <= NOT \ConfigureCodec|R.Data\(5);
\ConfigureCodec|ALT_INV_R.Data\(9) <= NOT \ConfigureCodec|R.Data\(9);
\ConfigureCodec|ALT_INV_R.Data\(1) <= NOT \ConfigureCodec|R.Data\(1);
\ConfigureCodec|ALT_INV_Mux9~1_combout\ <= NOT \ConfigureCodec|Mux9~1_combout\;
\ConfigureCodec|ALT_INV_R.Data\(14) <= NOT \ConfigureCodec|R.Data\(14);
\ConfigureCodec|ALT_INV_R.Data\(6) <= NOT \ConfigureCodec|R.Data\(6);
\ConfigureCodec|ALT_INV_R.Data\(10) <= NOT \ConfigureCodec|R.Data\(10);
\ConfigureCodec|ALT_INV_R.Data\(2) <= NOT \ConfigureCodec|R.Data\(2);
\ConfigureCodec|ALT_INV_Mux9~0_combout\ <= NOT \ConfigureCodec|Mux9~0_combout\;
\ConfigureCodec|ALT_INV_R.Data\(4) <= NOT \ConfigureCodec|R.Data\(4);
\ConfigureCodec|ALT_INV_R.Data\(0) <= NOT \ConfigureCodec|R.Data\(0);
\ConfigureCodec|ALT_INV_R.Data\(12) <= NOT \ConfigureCodec|R.Data\(12);
\TheI2sToPar|ALT_INV_LrcDlyd~q\ <= NOT \TheI2sToPar|LrcDlyd~q\;
\TheRxFsk|Lowpass|ALT_INV_R.SumState.Idle~q\ <= NOT \TheRxFsk|Lowpass|R.SumState.Idle~q\;
\TheRxFsk|Bandpasses:11:Bandpass0|ALT_INV_R.ValWet~q\ <= NOT \TheRxFsk|Bandpasses:11:Bandpass0|R.ValWet~q\;
\TheRxFsk|Lowpass|ALT_INV_R.SumState.SumEnable~q\ <= NOT \TheRxFsk|Lowpass|R.SumState.SumEnable~q\;
\TheRxFsk|Lowpass|ALT_INV_MultResultDelayed\(0) <= NOT \TheRxFsk|Lowpass|MultResultDelayed\(0);
\ConfigureCodec|ALT_INV_R.FrameState.Data1~q\ <= NOT \ConfigureCodec|R.FrameState.Data1~q\;
\ConfigureCodec|ALT_INV_NextR~9_combout\ <= NOT \ConfigureCodec|NextR~9_combout\;
\ConfigureCodec|ALT_INV_R.FrameState.RWBit~q\ <= NOT \ConfigureCodec|R.FrameState.RWBit~q\;
\ConfigureCodec|ALT_INV_NextR~8_combout\ <= NOT \ConfigureCodec|NextR~8_combout\;
\ConfigureCodec|ALT_INV_R.BitCtr\(0) <= NOT \ConfigureCodec|R.BitCtr\(0);
\ConfigureCodec|ALT_INV_R.BitCtr\(1) <= NOT \ConfigureCodec|R.BitCtr\(1);
\ConfigureCodec|ALT_INV_R.BitCtr\(2) <= NOT \ConfigureCodec|R.BitCtr\(2);
\ConfigureCodec|ALT_INV_R.BitCtr\(3) <= NOT \ConfigureCodec|R.BitCtr\(3);
\ConfigureCodec|ALT_INV_R.FrameState.Data2~q\ <= NOT \ConfigureCodec|R.FrameState.Data2~q\;
\ConfigureCodec|ALT_INV_R.Sdin~q\ <= NOT \ConfigureCodec|R.Sdin~q\;
\TheI2sToPar|ALT_INV_Decoder0~4_combout\ <= NOT \TheI2sToPar|Decoder0~4_combout\;
\TheI2sToPar|ALT_INV_D[14]~7_combout\ <= NOT \TheI2sToPar|D[14]~7_combout\;
\TheI2sToPar|ALT_INV_Decoder0~3_combout\ <= NOT \TheI2sToPar|Decoder0~3_combout\;
\TheI2sToPar|ALT_INV_Decoder0~2_combout\ <= NOT \TheI2sToPar|Decoder0~2_combout\;
\TheI2sToPar|ALT_INV_Decoder0~1_combout\ <= NOT \TheI2sToPar|Decoder0~1_combout\;
\TheI2sToPar|ALT_INV_Equal0~2_combout\ <= NOT \TheI2sToPar|Equal0~2_combout\;
\TheI2sToPar|ALT_INV_Equal0~1_combout\ <= NOT \TheI2sToPar|Equal0~1_combout\;
\TheI2sToPar|ALT_INV_BclkRiseEdge~combout\ <= NOT \TheI2sToPar|BclkRiseEdge~combout\;
\TheI2sToPar|ALT_INV_Equal0~0_combout\ <= NOT \TheI2sToPar|Equal0~0_combout\;
\TheI2sToPar|ALT_INV_AudioBitCtr\(0) <= NOT \TheI2sToPar|AudioBitCtr\(0);
\TheI2sToPar|ALT_INV_AudioBitCtr\(1) <= NOT \TheI2sToPar|AudioBitCtr\(1);
\TheI2sToPar|ALT_INV_AudioBitCtr\(2) <= NOT \TheI2sToPar|AudioBitCtr\(2);
\TheI2sToPar|ALT_INV_Decoder0~0_combout\ <= NOT \TheI2sToPar|Decoder0~0_combout\;
\TheI2sToPar|ALT_INV_State~q\ <= NOT \TheI2sToPar|State~q\;
\TheI2sToPar|ALT_INV_AudioBitCtr\(4) <= NOT \TheI2sToPar|AudioBitCtr\(4);
\TheI2sToPar|ALT_INV_AudioBitCtr\(3) <= NOT \TheI2sToPar|AudioBitCtr\(3);
\TheRxFsk|Lowpass|ALT_INV_R.EnableSumUp~q\ <= NOT \TheRxFsk|Lowpass|R.EnableSumUp~q\;
\TheRxFsk|Lowpass|ALT_INV_R.SelSumUp~q\ <= NOT \TheRxFsk|Lowpass|R.SelSumUp~q\;
\TheRxFsk|Lowpass|ALT_INV_R.SumState.SumWait2~q\ <= NOT \TheRxFsk|Lowpass|R.SumState.SumWait2~q\;
\TheRxFsk|Lowpass|ALT_INV_R.SumState.SumValid~q\ <= NOT \TheRxFsk|Lowpass|R.SumState.SumValid~q\;
\ConfigureCodec|ALT_INV_NextStateAndOutput:vSclkFalling~0_combout\ <= NOT \ConfigureCodec|NextStateAndOutput:vSclkFalling~0_combout\;
\ConfigureCodec|ALT_INV_Selector13~0_combout\ <= NOT \ConfigureCodec|Selector13~0_combout\;
\ConfigureCodec|ALT_INV_R.FrameState.Ack2~q\ <= NOT \ConfigureCodec|R.FrameState.Ack2~q\;
\ConfigureCodec|ALT_INV_R.FrameState.Ack1~q\ <= NOT \ConfigureCodec|R.FrameState.Ack1~q\;
\ConfigureCodec|ALT_INV_R.FrameState.Ack3~q\ <= NOT \ConfigureCodec|R.FrameState.Ack3~q\;
\ConfigureCodec|ALT_INV_R.Activity~0_combout\ <= NOT \ConfigureCodec|R.Activity~0_combout\;
\ConfigureCodec|ALT_INV_Selector16~0_combout\ <= NOT \ConfigureCodec|Selector16~0_combout\;
\GenStrobeI2C|ALT_INV_ClkCounter\(0) <= NOT \GenStrobeI2C|ClkCounter\(0);
\GenStrobeI2C|ALT_INV_ClkCounter\(1) <= NOT \GenStrobeI2C|ClkCounter\(1);
\GenStrobeI2C|ALT_INV_ClkCounter\(2) <= NOT \GenStrobeI2C|ClkCounter\(2);
\GenStrobeI2C|ALT_INV_ClkCounter\(3) <= NOT \GenStrobeI2C|ClkCounter\(3);
\GenStrobeI2C|ALT_INV_ClkCounter\(4) <= NOT \GenStrobeI2C|ClkCounter\(4);
\GenStrobeI2C|ALT_INV_ClkCounter\(5) <= NOT \GenStrobeI2C|ClkCounter\(5);
\GenClks|ALT_INV_Equal0~0_combout\ <= NOT \GenClks|Equal0~0_combout\;
\GenClks|ALT_INV_BitCounter\(3) <= NOT \GenClks|BitCounter\(3);
\GenClks|ALT_INV_BitCounter\(4) <= NOT \GenClks|BitCounter\(4);
\GenClks|ALT_INV_BitCounter\(5) <= NOT \GenClks|BitCounter\(5);
\GenClks|ALT_INV_BitCounter\(6) <= NOT \GenClks|BitCounter\(6);
\GenClks|ALT_INV_BitCounter\(7) <= NOT \GenClks|BitCounter\(7);
\GenClks|ALT_INV_BitCounter\(0) <= NOT \GenClks|BitCounter\(0);
\GenClks|ALT_INV_BitCounter\(1) <= NOT \GenClks|BitCounter\(1);
\GenClks|ALT_INV_BitCounter\(2) <= NOT \GenClks|BitCounter\(2);
\GenClks|ALT_INV_ADClrc~0_combout\ <= NOT \GenClks|ADClrc~0_combout\;
\TheParToI2s|ALT_INV_NextState~6_combout\ <= NOT \TheParToI2s|NextState~6_combout\;
\TheParToI2s|ALT_INV_Selector9~0_combout\ <= NOT \TheParToI2s|Selector9~0_combout\;
\TheParToI2s|ALT_INV_Selector7~0_combout\ <= NOT \TheParToI2s|Selector7~0_combout\;
\TheParToI2s|ALT_INV_Add0~0_combout\ <= NOT \TheParToI2s|Add0~0_combout\;
\TheI2sToPar|ALT_INV_D\(15) <= NOT \TheI2sToPar|D\(15);
\TheI2sToPar|ALT_INV_D\(7) <= NOT \TheI2sToPar|D\(7);
\TheI2sToPar|ALT_INV_D\(13) <= NOT \TheI2sToPar|D\(13);
\TheI2sToPar|ALT_INV_D\(5) <= NOT \TheI2sToPar|D\(5);
\TheI2sToPar|ALT_INV_D\(11) <= NOT \TheI2sToPar|D\(11);
\TheI2sToPar|ALT_INV_D\(3) <= NOT \TheI2sToPar|D\(3);
\TheI2sToPar|ALT_INV_D\(9) <= NOT \TheI2sToPar|D\(9);
\TheI2sToPar|ALT_INV_D\(1) <= NOT \TheI2sToPar|D\(1);
\TheI2sToPar|ALT_INV_D\(14) <= NOT \TheI2sToPar|D\(14);
\TheI2sToPar|ALT_INV_D\(6) <= NOT \TheI2sToPar|D\(6);
\TheI2sToPar|ALT_INV_D\(12) <= NOT \TheI2sToPar|D\(12);
\TheI2sToPar|ALT_INV_D\(4) <= NOT \TheI2sToPar|D\(4);
\TheParToI2s|ALT_INV_Selector8~0_combout\ <= NOT \TheParToI2s|Selector8~0_combout\;
\TheParToI2s|ALT_INV_NextBclkCtr~1_combout\ <= NOT \TheParToI2s|NextBclkCtr~1_combout\;
\TheParToI2s|ALT_INV_Selector6~1_combout\ <= NOT \TheParToI2s|Selector6~1_combout\;
\TheParToI2s|ALT_INV_NextBclkCtr~0_combout\ <= NOT \TheParToI2s|NextBclkCtr~0_combout\;
\TheParToI2s|ALT_INV_State.SyncingToBclk~q\ <= NOT \TheParToI2s|State.SyncingToBclk~q\;
\TheParToI2s|ALT_INV_State.WaitingValL~q\ <= NOT \TheParToI2s|State.WaitingValL~q\;
\TheParToI2s|ALT_INV_Selector6~0_combout\ <= NOT \TheParToI2s|Selector6~0_combout\;
\TheI2sToPar|ALT_INV_BclkDlyd~q\ <= NOT \TheI2sToPar|BclkDlyd~q\;
\TheParToI2s|ALT_INV_State.FirstBitEmptyR~q\ <= NOT \TheParToI2s|State.FirstBitEmptyR~q\;
\TheI2sToPar|ALT_INV_D\(10) <= NOT \TheI2sToPar|D\(10);
\TheI2sToPar|ALT_INV_D\(2) <= NOT \TheI2sToPar|D\(2);
\TheI2sToPar|ALT_INV_D\(8) <= NOT \TheI2sToPar|D\(8);
\TheI2sToPar|ALT_INV_ValL~q\ <= NOT \TheI2sToPar|ValL~q\;
\TheI2sToPar|ALT_INV_D\(0) <= NOT \TheI2sToPar|D\(0);
\GenClks|ALT_INV_ClkCounter\(0) <= NOT \GenClks|ClkCounter\(0);
\TheRxFsk|Lowpass|ALT_INV_R.ValWet~q\ <= NOT \TheRxFsk|Lowpass|R.ValWet~q\;
\ConfigureCodec|ALT_INV_R.AddrCtr[6]~1_combout\ <= NOT \ConfigureCodec|R.AddrCtr[6]~1_combout\;
\ConfigureCodec|ALT_INV_R.FrameState.Stop~q\ <= NOT \ConfigureCodec|R.FrameState.Stop~q\;
\ConfigureCodec|ALT_INV_R.AckError~q\ <= NOT \ConfigureCodec|R.AckError~q\;
\ConfigureCodec|ALT_INV_R.Sclk~q\ <= NOT \ConfigureCodec|R.Sclk~q\;
\ConfigureCodec|ALT_INV_Equal0~1_combout\ <= NOT \ConfigureCodec|Equal0~1_combout\;
\ConfigureCodec|ALT_INV_R.AddrCtr[6]~0_combout\ <= NOT \ConfigureCodec|R.AddrCtr[6]~0_combout\;
\ConfigureCodec|ALT_INV_R.FrameState.Idle~q\ <= NOT \ConfigureCodec|R.FrameState.Idle~q\;
\ConfigureCodec|ALT_INV_R.Activity~q\ <= NOT \ConfigureCodec|R.Activity~q\;
\ConfigureCodec|ALT_INV_Equal0~0_combout\ <= NOT \ConfigureCodec|Equal0~0_combout\;
ALT_INV_WaitCtr(0) <= NOT WaitCtr(0);
ALT_INV_WaitCtr(1) <= NOT WaitCtr(1);
\GenStrobeI2C|ALT_INV_oStrobe~q\ <= NOT \GenStrobeI2C|oStrobe~q\;
\TheParToI2s|ALT_INV_oLrc~0_combout\ <= NOT \TheParToI2s|oLrc~0_combout\;
\TheParToI2s|ALT_INV_State.FirstBitEmptyL~q\ <= NOT \TheParToI2s|State.FirstBitEmptyL~q\;
\GenClks|ALT_INV_ADClrc~q\ <= NOT \GenClks|ADClrc~q\;
\TheParToI2s|ALT_INV_Selector10~0_combout\ <= NOT \TheParToI2s|Selector10~0_combout\;
\TheParToI2s|ALT_INV_State.SendingR~q\ <= NOT \TheParToI2s|State.SendingR~q\;
\TheParToI2s|ALT_INV_State.SendingL~q\ <= NOT \TheParToI2s|State.SendingL~q\;
\TheParToI2s|ALT_INV_BclkCtr\(0) <= NOT \TheParToI2s|BclkCtr\(0);
\TheParToI2s|ALT_INV_BclkCtr\(2) <= NOT \TheParToI2s|BclkCtr\(2);
\TheParToI2s|ALT_INV_Mux1~3_combout\ <= NOT \TheParToI2s|Mux1~3_combout\;
\TheParToI2s|ALT_INV_LastValidDL\(15) <= NOT \TheParToI2s|LastValidDL\(15);
\TheParToI2s|ALT_INV_LastValidDL\(7) <= NOT \TheParToI2s|LastValidDL\(7);
\TheParToI2s|ALT_INV_LastValidDL\(13) <= NOT \TheParToI2s|LastValidDL\(13);
\TheParToI2s|ALT_INV_LastValidDL\(5) <= NOT \TheParToI2s|LastValidDL\(5);
\TheParToI2s|ALT_INV_Mux1~2_combout\ <= NOT \TheParToI2s|Mux1~2_combout\;
\TheParToI2s|ALT_INV_LastValidDL\(11) <= NOT \TheParToI2s|LastValidDL\(11);
\TheParToI2s|ALT_INV_LastValidDL\(3) <= NOT \TheParToI2s|LastValidDL\(3);
\TheParToI2s|ALT_INV_LastValidDL\(9) <= NOT \TheParToI2s|LastValidDL\(9);
\TheParToI2s|ALT_INV_LastValidDL\(1) <= NOT \TheParToI2s|LastValidDL\(1);
\TheParToI2s|ALT_INV_Mux1~1_combout\ <= NOT \TheParToI2s|Mux1~1_combout\;
\TheParToI2s|ALT_INV_LastValidDL\(14) <= NOT \TheParToI2s|LastValidDL\(14);
\TheParToI2s|ALT_INV_LastValidDL\(6) <= NOT \TheParToI2s|LastValidDL\(6);
\TheParToI2s|ALT_INV_LastValidDL\(12) <= NOT \TheParToI2s|LastValidDL\(12);
\TheParToI2s|ALT_INV_LastValidDL\(4) <= NOT \TheParToI2s|LastValidDL\(4);
\TheParToI2s|ALT_INV_Mux1~0_combout\ <= NOT \TheParToI2s|Mux1~0_combout\;
\TheParToI2s|ALT_INV_BclkCtr\(1) <= NOT \TheParToI2s|BclkCtr\(1);
\TheParToI2s|ALT_INV_BclkCtr\(3) <= NOT \TheParToI2s|BclkCtr\(3);
\TheParToI2s|ALT_INV_LastValidDL\(10) <= NOT \TheParToI2s|LastValidDL\(10);
\TheParToI2s|ALT_INV_LastValidDL\(2) <= NOT \TheParToI2s|LastValidDL\(2);
\TheParToI2s|ALT_INV_LastValidDL\(8) <= NOT \TheParToI2s|LastValidDL\(8);
\TheParToI2s|ALT_INV_LastValidDL\(0) <= NOT \TheParToI2s|LastValidDL\(0);
\GenClks|ALT_INV_BMclk~q\ <= NOT \GenClks|BMclk~q\;
\TheRxFsk|ALT_INV_oD~q\ <= NOT \TheRxFsk|oD~q\;
\ConfigureCodec|ALT_INV_R.Configured~q\ <= NOT \ConfigureCodec|R.Configured~q\;
\ALT_INV_Start~q\ <= NOT \Start~q\;
\SyncSwitchInput|ALT_INV_Metastable\(1) <= NOT \SyncSwitchInput|Metastable\(1);
\TheRxFsk|Lowpass|ALT_INV_Sum[-15]~q\ <= NOT \TheRxFsk|Lowpass|Sum[-15]~q\;
\TheRxFsk|Lowpass|ALT_INV_Sum[-14]~q\ <= NOT \TheRxFsk|Lowpass|Sum[-14]~q\;
\TheRxFsk|Lowpass|ALT_INV_Add4~61_sumout\ <= NOT \TheRxFsk|Lowpass|Add4~61_sumout\;
\TheRxFsk|Lowpass|ALT_INV_Sum[-13]~q\ <= NOT \TheRxFsk|Lowpass|Sum[-13]~q\;
\TheRxFsk|Lowpass|ALT_INV_Add4~57_sumout\ <= NOT \TheRxFsk|Lowpass|Add4~57_sumout\;
\TheRxFsk|Lowpass|ALT_INV_Sum[-12]~q\ <= NOT \TheRxFsk|Lowpass|Sum[-12]~q\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add0~33_sumout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Add0~33_sumout\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add0~5_sumout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Add0~5_sumout\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add1~33_sumout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Add1~33_sumout\;
\TheRxFsk|Lowpass|ALT_INV_Add4~53_sumout\ <= NOT \TheRxFsk|Lowpass|Add4~53_sumout\;
\TheRxFsk|Lowpass|ALT_INV_Sum[-11]~q\ <= NOT \TheRxFsk|Lowpass|Sum[-11]~q\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.WriteAddress\(7) <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(7);
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.WriteAddress\(6) <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(6);
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.WriteAddress\(5) <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(5);
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.WriteAddress\(4) <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(4);
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.WriteAddress\(3) <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(3);
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.WriteAddress\(2) <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(2);
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.WriteAddress\(1) <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(1);
\TheRxFsk|Lowpass|ALT_INV_Add4~49_sumout\ <= NOT \TheRxFsk|Lowpass|Add4~49_sumout\;
\TheRxFsk|Lowpass|ALT_INV_Sum[-10]~q\ <= NOT \TheRxFsk|Lowpass|Sum[-10]~q\;
\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a13\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a13\;
\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a14\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a14\;
\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a15\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a15\;
\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a1\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a1\;
\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a2\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a2\;
\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a3\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a3\;
\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a4\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a4\;
\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a5\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a5\;
\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a6\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a6\;
\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a7\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a7\;
\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a8\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a8\;
\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a9\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a9\;
\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a12~portbdataout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a12~portbdataout\;
\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a10\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a10\;
\TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a8\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a8\;
\TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a9\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a9\;
\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a11\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a11\;
\TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a10\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a10\;
\TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a11\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a11\;
\TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a12\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a12\;
\TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a13\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a13\;
\TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a14\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a14\;
\TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a15\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a15\;
\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a0~portbdataout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a0~portbdataout\;
\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a5\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a5\;
\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a6\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a6\;
\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a7\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a7\;
\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a8\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a8\;
\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a9\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a9\;
\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a10\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a10\;
\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a11\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a11\;
\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a12\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a12\;
\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a13\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a13\;
\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a14\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a14\;
\TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a0\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a0\;
\TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a1\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a1\;
\TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a2\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a2\;
\TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a3\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a3\;
\TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a4\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a4\;
\TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a5\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a5\;
\TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a6\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a6\;
\TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a7\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a7\;
\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a15\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a15\;
\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a1\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a1\;
\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a2\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a2\;
\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a3\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a3\;
\TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a0\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a0\;
\TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a1\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a1\;
\TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a2\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a2\;
\TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a3\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a3\;
\TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a4\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a4\;
\TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a5\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a5\;
\TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a6\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a6\;
\TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a7\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a7\;
\TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a8\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a8\;
\TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a9\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a9\;
\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a4~portbdataout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a4~portbdataout\;
\TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a10\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a10\;
\TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a11\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a11\;
\TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a12\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a12\;
\TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a13\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a13\;
\TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a14\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a14\;
\TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a15\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a15\;
\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a0~portbdataout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a0~portbdataout\;
\TheRxFsk|Lowpass|ALT_INV_Add4~45_sumout\ <= NOT \TheRxFsk|Lowpass|Add4~45_sumout\;
\TheRxFsk|Lowpass|ALT_INV_Sum[-9]~q\ <= NOT \TheRxFsk|Lowpass|Sum[-9]~q\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~39\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~39\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~38\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~38\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~37\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~37\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~36\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~36\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~35\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~35\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~34\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~34\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~33\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~33\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~32\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~32\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~31\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~31\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~30\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~30\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~29\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~29\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~28\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~28\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~27\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~27\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~26\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~26\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~25\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~25\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~24\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~24\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~23\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~23\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~22\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~22\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~21\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~21\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~20\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~20\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~19\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~19\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~18\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~18\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~17\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~17\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~16\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~16\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~15\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~15\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~14\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~14\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~13\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~13\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~12\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~12\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~11\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~11\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~10\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~10\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~9\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~9\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~8_resulta\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_resulta\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~39\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~39\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~38\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~38\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~37\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~37\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~36\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~36\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~35\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~35\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~34\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~34\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~33\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~33\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~32\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~32\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~31\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~31\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~30\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~30\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~29\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~29\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~28\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~28\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~27\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~27\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~26\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~26\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~25\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~25\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~24\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~24\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~23\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~23\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~22\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~22\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~21\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~21\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~20\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~20\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~19\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~19\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~18\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~18\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~17\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~17\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~16\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~16\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~15\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~15\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~14\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~14\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~13\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~13\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~12\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~12\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~11\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~11\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~10\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~10\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~9\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~9\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~8_resulta\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_resulta\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~39\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~39\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~38\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~38\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~37\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~37\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~36\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~36\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~35\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~35\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~34\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~34\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~33\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~33\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~32\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~32\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~31\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~31\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~30\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~30\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~29\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~29\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~28\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~28\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~27\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~27\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~26\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~26\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~25\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~25\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~24\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~24\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~23\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~23\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~22\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~22\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~21\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~21\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~20\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~20\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~19\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~19\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~18\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~18\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~17\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~17\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~16\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~16\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~15\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~15\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~14\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~14\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~13\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~13\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~12\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~12\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~11\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~11\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~10\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~10\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~9\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~9\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~8_resulta\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_resulta\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~39\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~39\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~38\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~38\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~37\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~37\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~36\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~36\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~35\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~35\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~34\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~34\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~33\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~33\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~32\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~32\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~31\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~31\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~30\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~30\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~29\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~29\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~28\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~28\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~27\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~27\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~26\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~26\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~25\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~25\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~24\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~24\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~23\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~23\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~22\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~22\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~21\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~21\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~20\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~20\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~19\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~19\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~18\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~18\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~17\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~17\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~16\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~16\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~15\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~15\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~14\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~14\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~13\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~13\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~12\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~12\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~11\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~11\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~10\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~10\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~9\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~9\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~8_resulta\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_resulta\;
\TheRxFsk|Lowpass|ALT_INV_Add4~41_sumout\ <= NOT \TheRxFsk|Lowpass|Add4~41_sumout\;
\TheRxFsk|Lowpass|ALT_INV_Sum[-8]~q\ <= NOT \TheRxFsk|Lowpass|Sum[-8]~q\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add3~1_sumout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Add3~1_sumout\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add3~1_sumout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Add3~1_sumout\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add3~1_sumout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Add3~1_sumout\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add3~1_sumout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Add3~1_sumout\;
\TheRxFsk|Lowpass|ALT_INV_Add4~37_sumout\ <= NOT \TheRxFsk|Lowpass|Add4~37_sumout\;
\TheRxFsk|Lowpass|ALT_INV_Sum[-7]~q\ <= NOT \TheRxFsk|Lowpass|Sum[-7]~q\;
\TheRxFsk|Lowpass|ALT_INV_Add4~33_sumout\ <= NOT \TheRxFsk|Lowpass|Add4~33_sumout\;
\TheRxFsk|Lowpass|ALT_INV_Sum[-6]~q\ <= NOT \TheRxFsk|Lowpass|Sum[-6]~q\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~65_sumout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Add4~65_sumout\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~65_sumout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Add4~65_sumout\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~65_sumout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Add4~65_sumout\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~65_sumout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Add4~65_sumout\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~61_sumout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Add4~61_sumout\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~61_sumout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Add4~61_sumout\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~61_sumout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Add4~61_sumout\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~61_sumout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Add4~61_sumout\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~57_sumout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Add4~57_sumout\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~57_sumout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Add4~57_sumout\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~57_sumout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Add4~57_sumout\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~57_sumout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Add4~57_sumout\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~53_sumout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Add4~53_sumout\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~53_sumout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Add4~53_sumout\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~53_sumout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Add4~53_sumout\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~53_sumout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Add4~53_sumout\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~49_sumout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Add4~49_sumout\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~49_sumout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Add4~49_sumout\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~49_sumout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Add4~49_sumout\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~49_sumout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Add4~49_sumout\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~45_sumout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Add4~45_sumout\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~45_sumout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Add4~45_sumout\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~45_sumout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Add4~45_sumout\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~45_sumout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Add4~45_sumout\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~41_sumout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Add4~41_sumout\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~41_sumout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Add4~41_sumout\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~41_sumout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Add4~41_sumout\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~41_sumout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Add4~41_sumout\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~37_sumout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Add4~37_sumout\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~37_sumout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Add4~37_sumout\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~37_sumout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Add4~37_sumout\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~37_sumout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Add4~37_sumout\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~33_sumout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Add4~33_sumout\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~33_sumout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Add4~33_sumout\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~33_sumout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Add4~33_sumout\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~33_sumout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Add4~33_sumout\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~29_sumout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Add4~29_sumout\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~29_sumout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Add4~29_sumout\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~29_sumout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Add4~29_sumout\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~29_sumout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Add4~29_sumout\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~25_sumout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Add4~25_sumout\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~25_sumout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Add4~25_sumout\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~25_sumout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Add4~25_sumout\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~25_sumout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Add4~25_sumout\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~21_sumout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Add4~21_sumout\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~21_sumout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Add4~21_sumout\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~21_sumout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Add4~21_sumout\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~21_sumout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Add4~21_sumout\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~17_sumout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Add4~17_sumout\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~17_sumout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Add4~17_sumout\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~17_sumout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Add4~17_sumout\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~17_sumout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Add4~17_sumout\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~13_sumout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Add4~13_sumout\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~13_sumout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Add4~13_sumout\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~13_sumout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Add4~13_sumout\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~13_sumout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Add4~13_sumout\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~5_sumout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Add4~5_sumout\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~5_sumout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Add4~5_sumout\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~1_sumout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Add4~1_sumout\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~1_sumout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Add4~1_sumout\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~5_sumout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Add4~5_sumout\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~5_sumout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Add4~5_sumout\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~1_sumout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Add4~1_sumout\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~1_sumout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Add4~1_sumout\;
\TheRxFsk|Lowpass|ALT_INV_Add4~29_sumout\ <= NOT \TheRxFsk|Lowpass|Add4~29_sumout\;
\TheRxFsk|Lowpass|ALT_INV_Sum[-5]~q\ <= NOT \TheRxFsk|Lowpass|Sum[-5]~q\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-1]~q\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-1]~q\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-1]~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-1]~q\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-1]~q\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-1]~q\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-1]~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-1]~q\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-2]~q\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-2]~q\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-2]~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-2]~q\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-2]~q\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-2]~q\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-2]~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-2]~q\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-3]~q\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-3]~q\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-3]~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-3]~q\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-3]~q\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-3]~q\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-3]~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-3]~q\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-4]~q\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-4]~q\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-4]~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-4]~q\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-4]~q\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-4]~q\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-4]~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-4]~q\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-5]~q\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-5]~q\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-5]~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-5]~q\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-5]~q\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-5]~q\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-5]~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-5]~q\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-6]~q\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-6]~q\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-6]~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-6]~q\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-6]~q\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-6]~q\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-6]~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-6]~q\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-7]~q\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-7]~q\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-7]~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-7]~q\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-7]~q\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-7]~q\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-7]~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-7]~q\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-8]~q\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-8]~q\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-8]~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-8]~q\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-8]~q\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-8]~q\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-8]~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-8]~q\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-9]~q\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-9]~q\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-9]~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-9]~q\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-9]~q\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-9]~q\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-9]~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-9]~q\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-10]~q\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-10]~q\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-10]~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-10]~q\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-10]~q\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-10]~q\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-10]~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-10]~q\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-11]~q\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-11]~q\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-11]~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-11]~q\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-11]~q\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-11]~q\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-11]~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-11]~q\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-12]~q\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-12]~q\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-12]~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-12]~q\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-12]~q\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-12]~q\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-12]~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-12]~q\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-13]~q\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-13]~q\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-13]~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-13]~q\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-13]~q\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-13]~q\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-13]~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-13]~q\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-14]~q\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-14]~q\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-14]~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-14]~q\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-14]~q\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-14]~q\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-14]~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-14]~q\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-15]~q\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-15]~q\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-15]~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-15]~q\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum\(0) <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Sum\(0);
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum\(0) <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Sum\(0);
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-15]~q\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-15]~q\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-15]~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-15]~q\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum\(0) <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|Sum\(0);
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum\(0) <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Sum\(0);
\TheRxFsk|Lowpass|ALT_INV_Add4~25_sumout\ <= NOT \TheRxFsk|Lowpass|Add4~25_sumout\;
\TheRxFsk|Lowpass|ALT_INV_Sum[-4]~q\ <= NOT \TheRxFsk|Lowpass|Sum[-4]~q\;
\TheRxFsk|ALT_INV_Add0~61_sumout\ <= NOT \TheRxFsk|Add0~61_sumout\;
\TheRxFsk|ALT_INV_Add1~61_sumout\ <= NOT \TheRxFsk|Add1~61_sumout\;
\TheRxFsk|ALT_INV_Add0~57_sumout\ <= NOT \TheRxFsk|Add0~57_sumout\;
\TheRxFsk|ALT_INV_Add1~57_sumout\ <= NOT \TheRxFsk|Add1~57_sumout\;
\TheRxFsk|ALT_INV_Add0~53_sumout\ <= NOT \TheRxFsk|Add0~53_sumout\;
\TheRxFsk|ALT_INV_Add1~53_sumout\ <= NOT \TheRxFsk|Add1~53_sumout\;
\TheRxFsk|ALT_INV_Add0~49_sumout\ <= NOT \TheRxFsk|Add0~49_sumout\;
\TheRxFsk|ALT_INV_Add1~49_sumout\ <= NOT \TheRxFsk|Add1~49_sumout\;
\TheRxFsk|ALT_INV_Add0~45_sumout\ <= NOT \TheRxFsk|Add0~45_sumout\;
\TheRxFsk|ALT_INV_Add1~45_sumout\ <= NOT \TheRxFsk|Add1~45_sumout\;
\TheRxFsk|ALT_INV_Add0~41_sumout\ <= NOT \TheRxFsk|Add0~41_sumout\;
\TheRxFsk|ALT_INV_Add1~41_sumout\ <= NOT \TheRxFsk|Add1~41_sumout\;
\TheRxFsk|ALT_INV_Add0~37_sumout\ <= NOT \TheRxFsk|Add0~37_sumout\;
\TheRxFsk|ALT_INV_Add1~37_sumout\ <= NOT \TheRxFsk|Add1~37_sumout\;
\TheRxFsk|ALT_INV_Add0~33_sumout\ <= NOT \TheRxFsk|Add0~33_sumout\;
\TheRxFsk|ALT_INV_Add1~33_sumout\ <= NOT \TheRxFsk|Add1~33_sumout\;
\TheRxFsk|ALT_INV_Add0~29_sumout\ <= NOT \TheRxFsk|Add0~29_sumout\;
\TheRxFsk|ALT_INV_Add1~29_sumout\ <= NOT \TheRxFsk|Add1~29_sumout\;
\TheRxFsk|ALT_INV_Add0~25_sumout\ <= NOT \TheRxFsk|Add0~25_sumout\;
\TheRxFsk|ALT_INV_Add1~25_sumout\ <= NOT \TheRxFsk|Add1~25_sumout\;
\TheRxFsk|ALT_INV_Add0~21_sumout\ <= NOT \TheRxFsk|Add0~21_sumout\;
\TheRxFsk|ALT_INV_Add1~21_sumout\ <= NOT \TheRxFsk|Add1~21_sumout\;
\TheRxFsk|ALT_INV_Add0~17_sumout\ <= NOT \TheRxFsk|Add0~17_sumout\;
\TheRxFsk|ALT_INV_Add1~17_sumout\ <= NOT \TheRxFsk|Add1~17_sumout\;
\TheRxFsk|ALT_INV_Add0~13_sumout\ <= NOT \TheRxFsk|Add0~13_sumout\;
\TheRxFsk|ALT_INV_Add1~13_sumout\ <= NOT \TheRxFsk|Add1~13_sumout\;
\TheRxFsk|ALT_INV_Add0~9_sumout\ <= NOT \TheRxFsk|Add0~9_sumout\;
\TheRxFsk|ALT_INV_Add1~9_sumout\ <= NOT \TheRxFsk|Add1~9_sumout\;
\TheRxFsk|Lowpass|ALT_INV_Add0~25_sumout\ <= NOT \TheRxFsk|Lowpass|Add0~25_sumout\;
\TheRxFsk|Lowpass|ALT_INV_Add0~13_sumout\ <= NOT \TheRxFsk|Lowpass|Add0~13_sumout\;
\TheRxFsk|Lowpass|ALT_INV_Add0~5_sumout\ <= NOT \TheRxFsk|Lowpass|Add0~5_sumout\;
\TheRxFsk|Lowpass|ALT_INV_Add1~25_sumout\ <= NOT \TheRxFsk|Lowpass|Add1~25_sumout\;
\TheRxFsk|Lowpass|ALT_INV_Add1~21_sumout\ <= NOT \TheRxFsk|Lowpass|Add1~21_sumout\;
\TheRxFsk|Lowpass|ALT_INV_Add1~17_sumout\ <= NOT \TheRxFsk|Lowpass|Add1~17_sumout\;
\TheRxFsk|Lowpass|ALT_INV_Add1~13_sumout\ <= NOT \TheRxFsk|Lowpass|Add1~13_sumout\;
\TheRxFsk|Lowpass|ALT_INV_Add1~9_sumout\ <= NOT \TheRxFsk|Lowpass|Add1~9_sumout\;
\TheRxFsk|Lowpass|ALT_INV_Add1~5_sumout\ <= NOT \TheRxFsk|Lowpass|Add1~5_sumout\;
\TheRxFsk|ALT_INV_Add0~5_sumout\ <= NOT \TheRxFsk|Add0~5_sumout\;
\TheRxFsk|ALT_INV_Add1~5_sumout\ <= NOT \TheRxFsk|Add1~5_sumout\;
\TheRxFsk|ALT_INV_Add0~1_sumout\ <= NOT \TheRxFsk|Add0~1_sumout\;
\TheRxFsk|ALT_INV_Add1~1_sumout\ <= NOT \TheRxFsk|Add1~1_sumout\;
\TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_Add2~29_sumout\ <= NOT \TheRxFsk|Bandpasses:0:Bandpass0|Add2~29_sumout\;
\TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_Add2~25_sumout\ <= NOT \TheRxFsk|Bandpasses:0:Bandpass0|Add2~25_sumout\;
\TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_Add2~21_sumout\ <= NOT \TheRxFsk|Bandpasses:0:Bandpass0|Add2~21_sumout\;
\TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_Add2~17_sumout\ <= NOT \TheRxFsk|Bandpasses:0:Bandpass0|Add2~17_sumout\;
\TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_Add2~13_sumout\ <= NOT \TheRxFsk|Bandpasses:0:Bandpass0|Add2~13_sumout\;
\TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_Add2~9_sumout\ <= NOT \TheRxFsk|Bandpasses:0:Bandpass0|Add2~9_sumout\;
\TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_Add2~5_sumout\ <= NOT \TheRxFsk|Bandpasses:0:Bandpass0|Add2~5_sumout\;
\TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_Add2~1_sumout\ <= NOT \TheRxFsk|Bandpasses:0:Bandpass0|Add2~1_sumout\;
\TheRxFsk|Lowpass|ALT_INV_Add4~21_sumout\ <= NOT \TheRxFsk|Lowpass|Add4~21_sumout\;
\TheRxFsk|Lowpass|ALT_INV_Sum[-3]~q\ <= NOT \TheRxFsk|Lowpass|Sum[-3]~q\;
\TheRxFsk|ALT_INV_Add2~65_sumout\ <= NOT \TheRxFsk|Add2~65_sumout\;
\TheRxFsk|ALT_INV_Add2~61_sumout\ <= NOT \TheRxFsk|Add2~61_sumout\;
\TheRxFsk|ALT_INV_Add2~57_sumout\ <= NOT \TheRxFsk|Add2~57_sumout\;
\TheRxFsk|ALT_INV_Add2~53_sumout\ <= NOT \TheRxFsk|Add2~53_sumout\;
\TheRxFsk|ALT_INV_Add2~49_sumout\ <= NOT \TheRxFsk|Add2~49_sumout\;
\TheRxFsk|ALT_INV_Add2~45_sumout\ <= NOT \TheRxFsk|Add2~45_sumout\;
\TheRxFsk|ALT_INV_Add2~41_sumout\ <= NOT \TheRxFsk|Add2~41_sumout\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[0]~DUPLICATE_q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[0]~DUPLICATE_q\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_R.SumState.Idle~DUPLICATE_q\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|R.SumState.Idle~DUPLICATE_q\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_R.SumState.SumEnable~DUPLICATE_q\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|R.SumState.SumEnable~DUPLICATE_q\;
\TheRxFsk|Lowpass|ALT_INV_R.ReadAddressSample[0]~DUPLICATE_q\ <= NOT \TheRxFsk|Lowpass|R.ReadAddressSample[0]~DUPLICATE_q\;
\TheRxFsk|Lowpass|ALT_INV_R.WriteAddress[1]~DUPLICATE_q\ <= NOT \TheRxFsk|Lowpass|R.WriteAddress[1]~DUPLICATE_q\;
\TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.ReadAddressCoef[0]~DUPLICATE_q\ <= NOT \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[0]~DUPLICATE_q\;
\TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.ReadAddressCoef[1]~DUPLICATE_q\ <= NOT \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[1]~DUPLICATE_q\;
\TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.ReadAddressCoef[2]~DUPLICATE_q\ <= NOT \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[2]~DUPLICATE_q\;
\TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.ReadAddressCoef[4]~DUPLICATE_q\ <= NOT \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[4]~DUPLICATE_q\;
\TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.ReadAddressCoef[5]~DUPLICATE_q\ <= NOT \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[5]~DUPLICATE_q\;
\TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.ReadAddressCoef[6]~DUPLICATE_q\ <= NOT \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[6]~DUPLICATE_q\;
\TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.ReadAddressCoef[7]~DUPLICATE_q\ <= NOT \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[7]~DUPLICATE_q\;
\TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef[6]~DUPLICATE_q\ <= NOT \TheRxFsk|Lowpass|R.ReadAddressCoef[6]~DUPLICATE_q\;
\ConfigureCodec|ALT_INV_R.FrameState.Data1~DUPLICATE_q\ <= NOT \ConfigureCodec|R.FrameState.Data1~DUPLICATE_q\;
\ConfigureCodec|ALT_INV_R.BitCtr[0]~DUPLICATE_q\ <= NOT \ConfigureCodec|R.BitCtr[0]~DUPLICATE_q\;
\ConfigureCodec|ALT_INV_R.BitCtr[3]~DUPLICATE_q\ <= NOT \ConfigureCodec|R.BitCtr[3]~DUPLICATE_q\;
\ConfigureCodec|ALT_INV_R.FrameState.Data2~DUPLICATE_q\ <= NOT \ConfigureCodec|R.FrameState.Data2~DUPLICATE_q\;
\TheI2sToPar|ALT_INV_AudioBitCtr[1]~DUPLICATE_q\ <= NOT \TheI2sToPar|AudioBitCtr[1]~DUPLICATE_q\;
\TheI2sToPar|ALT_INV_AudioBitCtr[2]~DUPLICATE_q\ <= NOT \TheI2sToPar|AudioBitCtr[2]~DUPLICATE_q\;
\TheRxFsk|Lowpass|ALT_INV_R.SumState.SumWait2~DUPLICATE_q\ <= NOT \TheRxFsk|Lowpass|R.SumState.SumWait2~DUPLICATE_q\;
\ConfigureCodec|ALT_INV_R.FrameState.Ack1~DUPLICATE_q\ <= NOT \ConfigureCodec|R.FrameState.Ack1~DUPLICATE_q\;
\GenStrobeI2C|ALT_INV_ClkCounter[0]~DUPLICATE_q\ <= NOT \GenStrobeI2C|ClkCounter[0]~DUPLICATE_q\;
\GenStrobeI2C|ALT_INV_ClkCounter[1]~DUPLICATE_q\ <= NOT \GenStrobeI2C|ClkCounter[1]~DUPLICATE_q\;
\GenClks|ALT_INV_BitCounter[1]~DUPLICATE_q\ <= NOT \GenClks|BitCounter[1]~DUPLICATE_q\;
\TheParToI2s|ALT_INV_State.SyncingToBclk~DUPLICATE_q\ <= NOT \TheParToI2s|State.SyncingToBclk~DUPLICATE_q\;
\ConfigureCodec|ALT_INV_R.FrameState.Idle~DUPLICATE_q\ <= NOT \ConfigureCodec|R.FrameState.Idle~DUPLICATE_q\;
\ALT_INV_WaitCtr[0]~DUPLICATE_q\ <= NOT \WaitCtr[0]~DUPLICATE_q\;
\TheParToI2s|ALT_INV_BclkCtr[2]~DUPLICATE_q\ <= NOT \TheParToI2s|BclkCtr[2]~DUPLICATE_q\;
\TheParToI2s|ALT_INV_BclkCtr[3]~DUPLICATE_q\ <= NOT \TheParToI2s|BclkCtr[3]~DUPLICATE_q\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-2]~DUPLICATE_q\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-2]~DUPLICATE_q\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-3]~DUPLICATE_q\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-3]~DUPLICATE_q\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-3]~DUPLICATE_q\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-3]~DUPLICATE_q\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-4]~DUPLICATE_q\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-4]~DUPLICATE_q\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-7]~DUPLICATE_q\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-7]~DUPLICATE_q\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-8]~DUPLICATE_q\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-8]~DUPLICATE_q\;
\ConfigureCodec|ALT_INV_R.AddrCtr[1]~DUPLICATE_q\ <= NOT \ConfigureCodec|R.AddrCtr[1]~DUPLICATE_q\;
\ConfigureCodec|ALT_INV_R.AddrCtr[2]~DUPLICATE_q\ <= NOT \ConfigureCodec|R.AddrCtr[2]~DUPLICATE_q\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-14]_OTERM179\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-14]_OTERM179\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-14]_OTERM177\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-14]_OTERM177\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-14]_OTERM175\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-14]_OTERM175\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-13]_OTERM173\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-13]_OTERM173\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-13]_OTERM171\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-13]_OTERM171\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-13]_OTERM169\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-13]_OTERM169\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-12]_OTERM167\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-12]_OTERM167\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-12]_OTERM165\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-12]_OTERM165\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-12]_OTERM163\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-12]_OTERM163\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-11]_OTERM161\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-11]_OTERM161\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-11]_OTERM159\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-11]_OTERM159\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-11]_OTERM157\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-11]_OTERM157\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-10]_OTERM155\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-10]_OTERM155\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-10]_OTERM153\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-10]_OTERM153\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-10]_OTERM151\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-10]_OTERM151\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-9]_OTERM149\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-9]_OTERM149\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-9]_OTERM147\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-9]_OTERM147\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-9]_OTERM145\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-9]_OTERM145\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-8]_OTERM143\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-8]_OTERM143\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-8]_OTERM141\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-8]_OTERM141\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-8]_OTERM139\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-8]_OTERM139\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-7]_OTERM137\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-7]_OTERM137\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-7]_OTERM135\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-7]_OTERM135\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-7]_OTERM133\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-7]_OTERM133\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-6]_OTERM131\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-6]_OTERM131\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-6]_OTERM129\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-6]_OTERM129\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-6]_OTERM127\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-6]_OTERM127\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-5]_OTERM125\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-5]_OTERM125\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-5]_OTERM123\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-5]_OTERM123\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-5]_OTERM121\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-5]_OTERM121\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-4]_OTERM119\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-4]_OTERM119\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-4]_OTERM117\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-4]_OTERM117\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-4]_OTERM115\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-4]_OTERM115\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-3]_OTERM113\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-3]_OTERM113\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-3]_OTERM111\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-3]_OTERM111\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-3]_OTERM109\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-3]_OTERM109\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-2]_OTERM107\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-2]_OTERM107\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-2]_OTERM105\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-2]_OTERM105\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-2]_OTERM103\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-2]_OTERM103\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-1]_OTERM101\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-1]_OTERM101\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-1]_OTERM99\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-1]_OTERM99\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-1]_OTERM97\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-1]_OTERM97\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-14]_OTERM95\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-14]_OTERM95\;
\TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-14]_OTERM93\ <= NOT \TheRxFsk|Lowpass|MultResultDelayed[-14]_OTERM93\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-13]_OTERM91\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-13]_OTERM91\;
\TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-13]_OTERM89\ <= NOT \TheRxFsk|Lowpass|MultResultDelayed[-13]_OTERM89\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM87\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM87\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM85\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM85\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM83\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM83\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM81\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM81\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM79\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM79\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM77\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM77\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM75\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM75\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM73\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM73\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM71\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM71\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM69\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM69\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM67\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM67\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM65\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM65\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-12]_OTERM63\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-12]_OTERM63\;
\TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-12]_OTERM61\ <= NOT \TheRxFsk|Lowpass|MultResultDelayed[-12]_OTERM61\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-11]_OTERM59\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-11]_OTERM59\;
\TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-11]_OTERM57\ <= NOT \TheRxFsk|Lowpass|MultResultDelayed[-11]_OTERM57\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-10]_OTERM55\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-10]_OTERM55\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-9]_OTERM53\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-9]_OTERM53\;
\TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-9]_OTERM51\ <= NOT \TheRxFsk|Lowpass|MultResultDelayed[-9]_OTERM51\;
\TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-10]_OTERM49\ <= NOT \TheRxFsk|Lowpass|MultResultDelayed[-10]_OTERM49\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-8]_OTERM47\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-8]_OTERM47\;
\TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-8]_OTERM45\ <= NOT \TheRxFsk|Lowpass|MultResultDelayed[-8]_OTERM45\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-7]_OTERM43\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-7]_OTERM43\;
\TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-7]_OTERM41\ <= NOT \TheRxFsk|Lowpass|MultResultDelayed[-7]_OTERM41\;
\TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-6]_OTERM39\ <= NOT \TheRxFsk|Lowpass|MultResultDelayed[-6]_OTERM39\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-6]_OTERM37\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-6]_OTERM37\;
\TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-5]_OTERM35\ <= NOT \TheRxFsk|Lowpass|MultResultDelayed[-5]_OTERM35\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-5]_OTERM33\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-5]_OTERM33\;
\TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-4]_OTERM31\ <= NOT \TheRxFsk|Lowpass|MultResultDelayed[-4]_OTERM31\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-4]_OTERM29\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-4]_OTERM29\;
\TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-3]_OTERM27\ <= NOT \TheRxFsk|Lowpass|MultResultDelayed[-3]_OTERM27\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-3]_OTERM25\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-3]_OTERM25\;
\TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-2]_OTERM23\ <= NOT \TheRxFsk|Lowpass|MultResultDelayed[-2]_OTERM23\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-2]_OTERM21\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-2]_OTERM21\;
\TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-1]_OTERM19\ <= NOT \TheRxFsk|Lowpass|MultResultDelayed[-1]_OTERM19\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-1]_OTERM17\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-1]_OTERM17\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM15\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM15\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM13\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM13\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM11\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM11\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM9\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM9\;
\TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM7\ <= NOT \TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM7\;
\TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM5\ <= NOT \TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM5\;
\TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM3\ <= NOT \TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM3\;
\TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM1\ <= NOT \TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM1\;
\ALT_INV_iADCdat~input_o\ <= NOT \iADCdat~input_o\;
\ALT_INV_inResetAsync~input_o\ <= NOT \inResetAsync~input_o\;
\ALT_INV_ioI2cSdin~input_o\ <= NOT \ioI2cSdin~input_o\;
\TheRxFsk|Lowpass|ALT_INV_CoefMemory~34_combout\ <= NOT \TheRxFsk|Lowpass|CoefMemory~34_combout\;
\TheRxFsk|Lowpass|ALT_INV_CoefMemory~33_combout\ <= NOT \TheRxFsk|Lowpass|CoefMemory~33_combout\;
\TheRxFsk|Lowpass|ALT_INV_CoefMemory~31_combout\ <= NOT \TheRxFsk|Lowpass|CoefMemory~31_combout\;
\TheRxFsk|Lowpass|ALT_INV_CoefMemory~30_combout\ <= NOT \TheRxFsk|Lowpass|CoefMemory~30_combout\;
\TheRxFsk|Lowpass|ALT_INV_CoefMemory~28_combout\ <= NOT \TheRxFsk|Lowpass|CoefMemory~28_combout\;
\TheRxFsk|Lowpass|ALT_INV_CoefMemory~27_combout\ <= NOT \TheRxFsk|Lowpass|CoefMemory~27_combout\;
\TheRxFsk|Lowpass|ALT_INV_CoefMemory~25_combout\ <= NOT \TheRxFsk|Lowpass|CoefMemory~25_combout\;
\TheRxFsk|Lowpass|ALT_INV_CoefMemory~24_combout\ <= NOT \TheRxFsk|Lowpass|CoefMemory~24_combout\;
\TheRxFsk|Lowpass|ALT_INV_CoefMemory~22_combout\ <= NOT \TheRxFsk|Lowpass|CoefMemory~22_combout\;
\TheRxFsk|Lowpass|ALT_INV_CoefMemory~21_combout\ <= NOT \TheRxFsk|Lowpass|CoefMemory~21_combout\;
\TheRxFsk|Lowpass|ALT_INV_CoefMemory~19_combout\ <= NOT \TheRxFsk|Lowpass|CoefMemory~19_combout\;
\TheRxFsk|Lowpass|ALT_INV_CoefMemory~18_combout\ <= NOT \TheRxFsk|Lowpass|CoefMemory~18_combout\;
\TheRxFsk|Lowpass|ALT_INV_CoefMemory~16_combout\ <= NOT \TheRxFsk|Lowpass|CoefMemory~16_combout\;
\TheRxFsk|Lowpass|ALT_INV_CoefMemory~15_combout\ <= NOT \TheRxFsk|Lowpass|CoefMemory~15_combout\;
\TheRxFsk|Lowpass|ALT_INV_CoefMemory~13_combout\ <= NOT \TheRxFsk|Lowpass|CoefMemory~13_combout\;
\TheRxFsk|Lowpass|ALT_INV_CoefMemory~12_combout\ <= NOT \TheRxFsk|Lowpass|CoefMemory~12_combout\;
\TheRxFsk|Lowpass|ALT_INV_CoefMemory~10_combout\ <= NOT \TheRxFsk|Lowpass|CoefMemory~10_combout\;
\TheRxFsk|Lowpass|ALT_INV_CoefMemory~9_combout\ <= NOT \TheRxFsk|Lowpass|CoefMemory~9_combout\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_vAdd~2_combout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|vAdd~2_combout\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_vAdd~1_combout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|vAdd~1_combout\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_vAdd~2_combout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|vAdd~2_combout\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_vAdd~1_combout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|vAdd~1_combout\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_vAdd~2_combout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|vAdd~2_combout\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_vAdd~1_combout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|vAdd~1_combout\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_vAdd~2_combout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|vAdd~2_combout\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_vAdd~1_combout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|vAdd~1_combout\;
\TheRxFsk|Lowpass|ALT_INV_vAdd~2_combout\ <= NOT \TheRxFsk|Lowpass|vAdd~2_combout\;
\TheRxFsk|Lowpass|ALT_INV_vAdd~1_combout\ <= NOT \TheRxFsk|Lowpass|vAdd~1_combout\;
\TheRxFsk|Lowpass|ALT_INV_vAdd~0_combout\ <= NOT \TheRxFsk|Lowpass|vAdd~0_combout\;
\TheRxFsk|Lowpass|ALT_INV_MultResult[-15]~14_combout\ <= NOT \TheRxFsk|Lowpass|MultResult[-15]~14_combout\;
\TheRxFsk|Lowpass|ALT_INV_MultResult[-14]~13_combout\ <= NOT \TheRxFsk|Lowpass|MultResult[-14]~13_combout\;
\TheRxFsk|Lowpass|ALT_INV_MultResult[-13]~12_combout\ <= NOT \TheRxFsk|Lowpass|MultResult[-13]~12_combout\;
\TheRxFsk|Lowpass|ALT_INV_MultResult[-12]~11_combout\ <= NOT \TheRxFsk|Lowpass|MultResult[-12]~11_combout\;
\TheRxFsk|Lowpass|ALT_INV_MultResult[-11]~10_combout\ <= NOT \TheRxFsk|Lowpass|MultResult[-11]~10_combout\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Equal0~0_combout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Equal0~0_combout\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Equal2~0_combout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|Equal2~0_combout\;
\TheRxFsk|Lowpass|ALT_INV_MultResult[-10]~9_combout\ <= NOT \TheRxFsk|Lowpass|MultResult[-10]~9_combout\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.ReadAddressSample\(8) <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(8);
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.ReadAddressSample\(7) <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(7);
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.ReadAddressSample\(6) <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(6);
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.ReadAddressSample\(5) <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(5);
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.ReadAddressSample\(4) <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(4);
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.ReadAddressSample\(3) <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(3);
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.ReadAddressSample\(2) <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(2);
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.ReadAddressSample\(1) <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(1);
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.ReadAddressSample\(0) <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(0);
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.WriteAddress\(8) <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(8);
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.WriteAddress\(0) <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(0);
\TheRxFsk|Lowpass|ALT_INV_MultResult[-9]~8_combout\ <= NOT \TheRxFsk|Lowpass|MultResult[-9]~8_combout\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed\(0) <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed\(0);
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-1]~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-1]~q\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-2]~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-2]~q\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-3]~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-3]~q\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-4]~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-4]~q\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-5]~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-5]~q\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-6]~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-6]~q\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-7]~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-7]~q\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-8]~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-8]~q\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-9]~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-9]~q\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-10]~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-10]~q\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-11]~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-11]~q\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-12]~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-12]~q\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-13]~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-13]~q\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-14]~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-14]~q\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-15]~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-15]~q\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\;
\TheRxFsk|Lowpass|ALT_INV_MultResult[-8]~7_combout\ <= NOT \TheRxFsk|Lowpass|MultResult[-8]~7_combout\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_vAdd~0_combout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|vAdd~0_combout\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_vAdd~0_combout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|vAdd~0_combout\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.SumState.SumSelect~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|R.SumState.SumSelect~q\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_R.SumState.SumSelect~q\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|R.SumState.SumSelect~q\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_vAdd~0_combout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|vAdd~0_combout\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_vAdd~0_combout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|vAdd~0_combout\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_R.SumState.SumSelect~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|R.SumState.SumSelect~q\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_R.SumState.SumSelect~q\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|R.SumState.SumSelect~q\;
\TheRxFsk|Lowpass|ALT_INV_MultResult[-7]~6_combout\ <= NOT \TheRxFsk|Lowpass|MultResult[-7]~6_combout\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResult[-1]~14_combout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-1]~14_combout\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResult[-1]~14_combout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-1]~14_combout\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResult[-1]~14_combout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-1]~14_combout\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResult[-1]~14_combout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-1]~14_combout\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResult[-2]~13_combout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-2]~13_combout\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResult[-2]~13_combout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-2]~13_combout\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResult[-2]~13_combout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-2]~13_combout\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResult[-2]~13_combout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-2]~13_combout\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResult[-3]~12_combout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-3]~12_combout\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResult[-3]~12_combout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-3]~12_combout\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResult[-3]~12_combout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-3]~12_combout\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResult[-3]~12_combout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-3]~12_combout\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResult[-4]~11_combout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-4]~11_combout\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResult[-4]~11_combout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-4]~11_combout\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResult[-4]~11_combout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-4]~11_combout\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResult[-4]~11_combout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-4]~11_combout\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResult[-5]~10_combout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-5]~10_combout\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResult[-5]~10_combout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-5]~10_combout\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResult[-5]~10_combout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-5]~10_combout\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResult[-5]~10_combout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-5]~10_combout\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResult[-6]~9_combout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-6]~9_combout\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResult[-6]~9_combout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-6]~9_combout\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResult[-6]~9_combout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-6]~9_combout\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResult[-6]~9_combout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-6]~9_combout\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResult[-7]~8_combout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-7]~8_combout\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResult[-7]~8_combout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-7]~8_combout\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResult[-7]~8_combout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-7]~8_combout\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResult[-7]~8_combout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-7]~8_combout\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResult[-8]~7_combout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-8]~7_combout\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResult[-8]~7_combout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-8]~7_combout\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResult[-8]~7_combout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-8]~7_combout\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResult[-8]~7_combout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-8]~7_combout\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResult[-9]~6_combout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-9]~6_combout\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResult[-9]~6_combout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-9]~6_combout\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResult[-9]~6_combout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-9]~6_combout\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResult[-9]~6_combout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-9]~6_combout\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResult[-10]~5_combout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-10]~5_combout\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResult[-10]~5_combout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-10]~5_combout\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResult[-10]~5_combout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-10]~5_combout\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResult[-10]~5_combout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-10]~5_combout\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResult[-11]~4_combout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-11]~4_combout\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResult[-11]~4_combout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-11]~4_combout\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResult[-11]~4_combout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-11]~4_combout\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResult[-11]~4_combout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-11]~4_combout\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResult[-12]~3_combout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-12]~3_combout\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResult[-12]~3_combout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-12]~3_combout\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResult[-12]~3_combout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-12]~3_combout\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResult[-12]~3_combout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-12]~3_combout\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResult[-13]~2_combout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-13]~2_combout\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResult[-13]~2_combout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-13]~2_combout\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResult[-13]~2_combout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-13]~2_combout\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResult[-13]~2_combout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-13]~2_combout\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResult[-14]~1_combout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-14]~1_combout\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResult[-14]~1_combout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-14]~1_combout\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResult[-14]~1_combout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-14]~1_combout\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResult[-14]~1_combout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-14]~1_combout\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResult[-15]~0_combout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-15]~0_combout\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResult[-15]~0_combout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-15]~0_combout\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.SumState.SumValid~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|R.SumState.SumValid~q\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_R.SumState.SumValid~q\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|R.SumState.SumValid~q\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResult[-15]~0_combout\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-15]~0_combout\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResult[-15]~0_combout\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-15]~0_combout\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_R.SumState.SumValid~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|R.SumState.SumValid~q\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_R.SumState.SumValid~q\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|R.SumState.SumValid~q\;
\TheRxFsk|Lowpass|ALT_INV_MultResult[-6]~5_combout\ <= NOT \TheRxFsk|Lowpass|MultResult[-6]~5_combout\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.SumState.Idle~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|R.SumState.Idle~q\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.SumState.SumEnable~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|R.SumState.SumEnable~q\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.SumState.SumWait2~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|R.SumState.SumWait2~q\;
\TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed\(0) <= NOT \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed\(0);
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_R.SumState.Idle~q\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|R.SumState.Idle~q\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_R.SumState.SumEnable~q\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|R.SumState.SumEnable~q\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_R.SumState.SumWait2~q\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|R.SumState.SumWait2~q\;
\TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed\(0) <= NOT \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed\(0);
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_R.SumState.Idle~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|R.SumState.Idle~q\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_R.SumState.SumEnable~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|R.SumState.SumEnable~q\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_R.SumState.SumWait2~q\ <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|R.SumState.SumWait2~q\;
\TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed\(0) <= NOT \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed\(0);
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_R.SumState.Idle~q\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|R.SumState.Idle~q\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_R.SumState.SumEnable~q\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|R.SumState.SumEnable~q\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_R.SumState.SumWait2~q\ <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|R.SumState.SumWait2~q\;
\TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed\(0) <= NOT \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed\(0);
\TheRxFsk|Lowpass|ALT_INV_MultResult[-5]~4_combout\ <= NOT \TheRxFsk|Lowpass|MultResult[-5]~4_combout\;

-- Location: IOOBUF_X12_Y81_N19
\oI2cSclk~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "true",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \ConfigureCodec|ALT_INV_R.Sclk~q\,
	devoe => ww_devoe,
	o => ww_oI2cSclk);

-- Location: IOOBUF_X89_Y8_N39
\oSEG0[0]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \SyncSwitchInput|Metastable\(1),
	devoe => ww_devoe,
	o => ww_oSEG0(0));

-- Location: IOOBUF_X89_Y11_N79
\oSEG0[1]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => GND,
	devoe => ww_devoe,
	o => ww_oSEG0(1));

-- Location: IOOBUF_X89_Y11_N96
\oSEG0[2]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => GND,
	devoe => ww_devoe,
	o => ww_oSEG0(2));

-- Location: IOOBUF_X89_Y4_N79
\oSEG0[3]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => VCC,
	devoe => ww_devoe,
	o => ww_oSEG0(3));

-- Location: IOOBUF_X89_Y13_N56
\oSEG0[4]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => VCC,
	devoe => ww_devoe,
	o => ww_oSEG0(4));

-- Location: IOOBUF_X89_Y13_N39
\oSEG0[5]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \SyncSwitchInput|ALT_INV_Metastable\(1),
	devoe => ww_devoe,
	o => ww_oSEG0(5));

-- Location: IOOBUF_X89_Y4_N96
\oSEG0[6]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \SyncSwitchInput|ALT_INV_Metastable\(1),
	devoe => ww_devoe,
	o => ww_oSEG0(6));

-- Location: IOOBUF_X89_Y6_N39
\oSEG1[0]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => GND,
	devoe => ww_devoe,
	o => ww_oSEG1(0));

-- Location: IOOBUF_X89_Y6_N56
\oSEG1[1]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => GND,
	devoe => ww_devoe,
	o => ww_oSEG1(1));

-- Location: IOOBUF_X89_Y16_N39
\oSEG1[2]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => GND,
	devoe => ww_devoe,
	o => ww_oSEG1(2));

-- Location: IOOBUF_X89_Y16_N56
\oSEG1[3]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => GND,
	devoe => ww_devoe,
	o => ww_oSEG1(3));

-- Location: IOOBUF_X89_Y15_N39
\oSEG1[4]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => GND,
	devoe => ww_devoe,
	o => ww_oSEG1(4));

-- Location: IOOBUF_X89_Y15_N56
\oSEG1[5]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => GND,
	devoe => ww_devoe,
	o => ww_oSEG1(5));

-- Location: IOOBUF_X89_Y8_N56
\oSEG1[6]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => VCC,
	devoe => ww_devoe,
	o => ww_oSEG1(6));

-- Location: IOOBUF_X89_Y9_N22
\oSEG2[0]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => GND,
	devoe => ww_devoe,
	o => ww_oSEG2(0));

-- Location: IOOBUF_X89_Y23_N39
\oSEG2[1]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => GND,
	devoe => ww_devoe,
	o => ww_oSEG2(1));

-- Location: IOOBUF_X89_Y23_N56
\oSEG2[2]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => GND,
	devoe => ww_devoe,
	o => ww_oSEG2(2));

-- Location: IOOBUF_X89_Y20_N79
\oSEG2[3]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => GND,
	devoe => ww_devoe,
	o => ww_oSEG2(3));

-- Location: IOOBUF_X89_Y25_N39
\oSEG2[4]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => GND,
	devoe => ww_devoe,
	o => ww_oSEG2(4));

-- Location: IOOBUF_X89_Y20_N96
\oSEG2[5]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => GND,
	devoe => ww_devoe,
	o => ww_oSEG2(5));

-- Location: IOOBUF_X89_Y25_N56
\oSEG2[6]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => VCC,
	devoe => ww_devoe,
	o => ww_oSEG2(6));

-- Location: IOOBUF_X89_Y16_N5
\oSEG3[0]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => GND,
	devoe => ww_devoe,
	o => ww_oSEG3(0));

-- Location: IOOBUF_X89_Y16_N22
\oSEG3[1]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => GND,
	devoe => ww_devoe,
	o => ww_oSEG3(1));

-- Location: IOOBUF_X89_Y4_N45
\oSEG3[2]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => GND,
	devoe => ww_devoe,
	o => ww_oSEG3(2));

-- Location: IOOBUF_X89_Y4_N62
\oSEG3[3]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => GND,
	devoe => ww_devoe,
	o => ww_oSEG3(3));

-- Location: IOOBUF_X89_Y21_N39
\oSEG3[4]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => GND,
	devoe => ww_devoe,
	o => ww_oSEG3(4));

-- Location: IOOBUF_X89_Y11_N62
\oSEG3[5]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => GND,
	devoe => ww_devoe,
	o => ww_oSEG3(5));

-- Location: IOOBUF_X89_Y9_N5
\oSEG3[6]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => VCC,
	devoe => ww_devoe,
	o => ww_oSEG3(6));

-- Location: IOOBUF_X89_Y11_N45
\oSEG4[0]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => GND,
	devoe => ww_devoe,
	o => ww_oSEG4(0));

-- Location: IOOBUF_X89_Y13_N5
\oSEG4[1]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => GND,
	devoe => ww_devoe,
	o => ww_oSEG4(1));

-- Location: IOOBUF_X89_Y13_N22
\oSEG4[2]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => GND,
	devoe => ww_devoe,
	o => ww_oSEG4(2));

-- Location: IOOBUF_X89_Y8_N22
\oSEG4[3]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => GND,
	devoe => ww_devoe,
	o => ww_oSEG4(3));

-- Location: IOOBUF_X89_Y15_N22
\oSEG4[4]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => GND,
	devoe => ww_devoe,
	o => ww_oSEG4(4));

-- Location: IOOBUF_X89_Y15_N5
\oSEG4[5]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => GND,
	devoe => ww_devoe,
	o => ww_oSEG4(5));

-- Location: IOOBUF_X89_Y20_N45
\oSEG4[6]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => VCC,
	devoe => ww_devoe,
	o => ww_oSEG4(6));

-- Location: IOOBUF_X89_Y20_N62
\oSEG5[0]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => GND,
	devoe => ww_devoe,
	o => ww_oSEG5(0));

-- Location: IOOBUF_X89_Y21_N56
\oSEG5[1]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => GND,
	devoe => ww_devoe,
	o => ww_oSEG5(1));

-- Location: IOOBUF_X89_Y25_N22
\oSEG5[2]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => GND,
	devoe => ww_devoe,
	o => ww_oSEG5(2));

-- Location: IOOBUF_X89_Y23_N22
\oSEG5[3]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => GND,
	devoe => ww_devoe,
	o => ww_oSEG5(3));

-- Location: IOOBUF_X89_Y9_N56
\oSEG5[4]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => GND,
	devoe => ww_devoe,
	o => ww_oSEG5(4));

-- Location: IOOBUF_X89_Y23_N5
\oSEG5[5]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => GND,
	devoe => ww_devoe,
	o => ww_oSEG5(5));

-- Location: IOOBUF_X89_Y9_N39
\oSEG5[6]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => VCC,
	devoe => ww_devoe,
	o => ww_oSEG5(6));

-- Location: IOOBUF_X52_Y0_N2
\oLed[0]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|locked_wire\(0),
	devoe => ww_devoe,
	o => ww_oLed(0));

-- Location: IOOBUF_X52_Y0_N19
\oLed[1]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \Start~q\,
	devoe => ww_devoe,
	o => ww_oLed(1));

-- Location: IOOBUF_X60_Y0_N2
\oLed[2]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \ConfigureCodec|R.Configured~DUPLICATE_q\,
	devoe => ww_devoe,
	o => ww_oLed(2));

-- Location: IOOBUF_X80_Y0_N2
\oLed[3]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \SyncSwitchInput|Metastable\(1),
	devoe => ww_devoe,
	o => ww_oLed(3));

-- Location: IOOBUF_X60_Y0_N19
\oLed[4]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \SyncSwitchInput|Metastable\(1),
	devoe => ww_devoe,
	o => ww_oLed(4));

-- Location: IOOBUF_X80_Y0_N19
\oLed[5]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \TheRxFsk|oD~q\,
	devoe => ww_devoe,
	o => ww_oLed(5));

-- Location: IOOBUF_X84_Y0_N2
\oLed[6]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => GND,
	devoe => ww_devoe,
	o => ww_oLed(6));

-- Location: IOOBUF_X89_Y6_N5
\oLed[7]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => GND,
	devoe => ww_devoe,
	o => ww_oLed(7));

-- Location: IOOBUF_X89_Y8_N5
\oLed[8]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => GND,
	devoe => ww_devoe,
	o => ww_oLed(8));

-- Location: IOOBUF_X89_Y6_N22
\oLed[9]~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => GND,
	devoe => ww_devoe,
	o => ww_oLed(9));

-- Location: IOOBUF_X2_Y81_N76
\oMclk~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \GenClks|BMclk~q\,
	devoe => ww_devoe,
	o => ww_oMclk);

-- Location: IOOBUF_X16_Y81_N19
\oBclk~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \GenClks|BMclk~q\,
	devoe => ww_devoe,
	o => ww_oBclk);

-- Location: IOOBUF_X16_Y81_N2
\oDACdat~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \TheParToI2s|Selector10~1_combout\,
	devoe => ww_devoe,
	o => ww_oDACdat);

-- Location: IOOBUF_X8_Y81_N19
\oADClrc~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \GenClks|ADClrc~q\,
	devoe => ww_devoe,
	o => ww_oADClrc);

-- Location: IOOBUF_X24_Y81_N2
\oDAClrc~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "false",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \TheParToI2s|ALT_INV_oLrc~0_combout\,
	devoe => ww_devoe,
	o => ww_oDAClrc);

-- Location: IOOBUF_X12_Y81_N2
\ioI2cSdin~output\ : cyclonev_io_obuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	open_drain_output => "true",
	shift_series_termination_control => "false")
-- pragma translate_on
PORT MAP (
	i => \ConfigureCodec|ALT_INV_R.Sdin~q\,
	oe => VCC,
	devoe => ww_devoe,
	o => ioI2cSdin);

-- Location: IOIBUF_X32_Y0_N1
\iClk~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_iClk,
	o => \iClk~input_o\);

-- Location: PLLREFCLKSELECT_X0_Y21_N0
\PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~PLL_REFCLK_SELECT\ : cyclonev_pll_refclk_select
-- pragma translate_off
GENERIC MAP (
	pll_auto_clk_sw_en => "false",
	pll_clk_loss_edge => "both_edges",
	pll_clk_loss_sw_en => "false",
	pll_clk_sw_dly => 0,
	pll_clkin_0_src => "clk_0",
	pll_clkin_1_src => "ref_clk1",
	pll_manu_clk_sw_en => "false",
	pll_sw_refclk_src => "clk_0")
-- pragma translate_on
PORT MAP (
	clkin => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~PLL_REFCLK_SELECT_CLKIN_bus\,
	clkout => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~PLL_REFCLK_SELECT_O_CLKOUT\,
	extswitchbuf => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~PLL_REFCLK_SELECT_O_EXTSWITCHBUF\);

-- Location: IOIBUF_X36_Y0_N1
\inResetAsync~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_inResetAsync,
	o => \inResetAsync~input_o\);

-- Location: FRACTIONALPLL_X0_Y15_N0
\PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL\ : cyclonev_fractional_pll
-- pragma translate_off
GENERIC MAP (
	dsm_accumulator_reset_value => 0,
	forcelock => "false",
	mimic_fbclk_type => "none",
	nreset_invert => "true",
	output_clock_frequency => "480.0 mhz",
	pll_atb => 0,
	pll_bwctrl => 10000,
	pll_cmp_buf_dly => "0 ps",
	pll_cp_comp => "true",
	pll_cp_current => 20,
	pll_ctrl_override_setting => "false",
	pll_dsm_dither => "disable",
	pll_dsm_out_sel => "disable",
	pll_dsm_reset => "false",
	pll_ecn_bypass => "false",
	pll_ecn_test_en => "false",
	pll_enable => "true",
	pll_fbclk_mux_1 => "glb",
	pll_fbclk_mux_2 => "m_cnt",
	pll_fractional_carry_out => 32,
	pll_fractional_division => 1,
	pll_fractional_division_string => "'0'",
	pll_fractional_value_ready => "true",
	pll_lf_testen => "false",
	pll_lock_fltr_cfg => 25,
	pll_lock_fltr_test => "false",
	pll_m_cnt_bypass_en => "false",
	pll_m_cnt_coarse_dly => "0 ps",
	pll_m_cnt_fine_dly => "0 ps",
	pll_m_cnt_hi_div => 24,
	pll_m_cnt_in_src => "ph_mux_clk",
	pll_m_cnt_lo_div => 24,
	pll_m_cnt_odd_div_duty_en => "false",
	pll_m_cnt_ph_mux_prst => 6,
	pll_m_cnt_prst => 5,
	pll_n_cnt_bypass_en => "false",
	pll_n_cnt_coarse_dly => "0 ps",
	pll_n_cnt_fine_dly => "0 ps",
	pll_n_cnt_hi_div => 3,
	pll_n_cnt_lo_div => 2,
	pll_n_cnt_odd_div_duty_en => "false",
	pll_ref_buf_dly => "0 ps",
	pll_reg_boost => 0,
	pll_regulator_bypass => "false",
	pll_ripplecap_ctrl => 0,
	pll_slf_rst => "false",
	pll_tclk_mux_en => "false",
	pll_tclk_sel => "n_src",
	pll_test_enable => "false",
	pll_testdn_enable => "false",
	pll_testup_enable => "false",
	pll_unlock_fltr_cfg => 2,
	pll_vco_div => 2,
	pll_vco_ph0_en => "true",
	pll_vco_ph1_en => "true",
	pll_vco_ph2_en => "true",
	pll_vco_ph3_en => "true",
	pll_vco_ph4_en => "true",
	pll_vco_ph5_en => "true",
	pll_vco_ph6_en => "true",
	pll_vco_ph7_en => "true",
	pll_vctrl_test_voltage => 750,
	reference_clock_frequency => "50.0 mhz",
	vccd0g_atb => "disable",
	vccd0g_output => 0,
	vccd1g_atb => "disable",
	vccd1g_output => 0,
	vccm1g_tap => 2,
	vccr_pd => "false",
	vcodiv_override => "false",
  fractional_pll_index => 0)
-- pragma translate_on
PORT MAP (
	coreclkfb => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|fboutclk_wire\(0),
	ecnc1test => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~PLL_REFCLK_SELECT_O_EXTSWITCHBUF\,
	nresync => \ALT_INV_inResetAsync~input_o\,
	refclkin => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~PLL_REFCLK_SELECT_O_CLKOUT\,
	shift => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~PLL_RECONFIG_O_SHIFT\,
	shiftdonein => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~PLL_RECONFIG_O_SHIFT\,
	shiften => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~PLL_RECONFIG_O_SHIFTENM\,
	up => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~PLL_RECONFIG_O_UP\,
	cntnen => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_CNTNEN\,
	fbclk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|fboutclk_wire\(0),
	lock => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|locked_wire\(0),
	tclk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_TCLK\,
	vcoph => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_VCOPH_bus\,
	mhi => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_MHI_bus\);

-- Location: PLLRECONFIG_X0_Y19_N0
\PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~PLL_RECONFIG\ : cyclonev_pll_reconfig
-- pragma translate_off
GENERIC MAP (
  fractional_pll_index => 0)
-- pragma translate_on
PORT MAP (
	cntnen => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_CNTNEN\,
	mhi => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~PLL_RECONFIG_MHI_bus\,
	shift => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~PLL_RECONFIG_O_SHIFT\,
	shiftenm => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~PLL_RECONFIG_O_SHIFTENM\,
	up => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~PLL_RECONFIG_O_UP\,
	shiften => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~PLL_RECONFIG_SHIFTEN_bus\);

-- Location: PLLOUTPUTCOUNTER_X0_Y20_N1
\PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~PLL_OUTPUT_COUNTER\ : cyclonev_pll_output_counter
-- pragma translate_off
GENERIC MAP (
	c_cnt_coarse_dly => "0 ps",
	c_cnt_fine_dly => "0 ps",
	c_cnt_in_src => "ph_mux_clk",
	c_cnt_ph_mux_prst => 0,
	c_cnt_prst => 1,
	cnt_fpll_src => "fpll_0",
	dprio0_cnt_bypass_en => "false",
	dprio0_cnt_hi_div => 5,
	dprio0_cnt_lo_div => 5,
	dprio0_cnt_odd_div_even_duty_en => "false",
	duty_cycle => 50,
	output_clock_frequency => "48.0 mhz",
	phase_shift => "0 ps",
  fractional_pll_index => 0,
  output_counter_index => 6)
-- pragma translate_on
PORT MAP (
	nen0 => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_CNTNEN\,
	shift0 => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~PLL_RECONFIG_O_SHIFT\,
	shiften => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~PLL_RECONFIGSHIFTEN6\,
	tclk0 => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~FRACTIONAL_PLL_O_TCLK\,
	up0 => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~PLL_RECONFIG_O_UP\,
	vco0ph => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|general[0].gpll~PLL_OUTPUT_COUNTER_VCO0PH_bus\,
	divclk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire\(0));

-- Location: CLKCTRL_G0
\PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0\ : cyclonev_clkena
-- pragma translate_off
GENERIC MAP (
	clock_type => "global clock",
	disable_mode => "low",
	ena_register_mode => "always enabled",
	ena_register_power_up => "high",
	test_syn => "high")
-- pragma translate_on
PORT MAP (
	inclk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire\(0),
	outclk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\);

-- Location: CLKCTRL_G6
\inResetAsync~inputCLKENA0\ : cyclonev_clkena
-- pragma translate_off
GENERIC MAP (
	clock_type => "global clock",
	disable_mode => "low",
	ena_register_mode => "always enabled",
	ena_register_power_up => "high",
	test_syn => "high")
-- pragma translate_on
PORT MAP (
	inclk => \inResetAsync~input_o\,
	outclk => \inResetAsync~inputCLKENA0_outclk\);

-- Location: FF_X18_Y66_N35
\GenStrobeI2C|ClkCounter[1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \GenStrobeI2C|ClkCounter[1]~4_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \GenStrobeI2C|ClkCounter\(1));

-- Location: FF_X18_Y66_N26
\GenStrobeI2C|ClkCounter[0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \GenStrobeI2C|ClkCounter[0]~5_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \GenStrobeI2C|ClkCounter\(0));

-- Location: LABCELL_X18_Y66_N24
\GenStrobeI2C|ClkCounter[0]~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \GenStrobeI2C|ClkCounter[0]~5_combout\ = ( !\GenStrobeI2C|ClkCounter\(0) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111111111111000000000000000011111111111111110000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datae => \GenStrobeI2C|ALT_INV_ClkCounter\(0),
	combout => \GenStrobeI2C|ClkCounter[0]~5_combout\);

-- Location: FF_X18_Y66_N25
\GenStrobeI2C|ClkCounter[0]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \GenStrobeI2C|ClkCounter[0]~5_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \GenStrobeI2C|ClkCounter[0]~DUPLICATE_q\);

-- Location: LABCELL_X18_Y66_N33
\GenStrobeI2C|ClkCounter[1]~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \GenStrobeI2C|ClkCounter[1]~4_combout\ = ( !\GenStrobeI2C|ClkCounter\(1) & ( \GenStrobeI2C|ClkCounter[0]~DUPLICATE_q\ ) ) # ( \GenStrobeI2C|ClkCounter\(1) & ( !\GenStrobeI2C|ClkCounter[0]~DUPLICATE_q\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111111111111111111110000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datae => \GenStrobeI2C|ALT_INV_ClkCounter\(1),
	dataf => \GenStrobeI2C|ALT_INV_ClkCounter[0]~DUPLICATE_q\,
	combout => \GenStrobeI2C|ClkCounter[1]~4_combout\);

-- Location: FF_X18_Y66_N34
\GenStrobeI2C|ClkCounter[1]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \GenStrobeI2C|ClkCounter[1]~4_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \GenStrobeI2C|ClkCounter[1]~DUPLICATE_q\);

-- Location: LABCELL_X18_Y66_N0
\GenStrobeI2C|ClkCounter[2]~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \GenStrobeI2C|ClkCounter[2]~3_combout\ = ( \GenStrobeI2C|ClkCounter\(2) & ( \GenStrobeI2C|ClkCounter[1]~DUPLICATE_q\ & ( !\GenStrobeI2C|ClkCounter\(0) ) ) ) # ( !\GenStrobeI2C|ClkCounter\(2) & ( \GenStrobeI2C|ClkCounter[1]~DUPLICATE_q\ & ( 
-- \GenStrobeI2C|ClkCounter\(0) ) ) ) # ( \GenStrobeI2C|ClkCounter\(2) & ( !\GenStrobeI2C|ClkCounter[1]~DUPLICATE_q\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100001111000011111111000011110000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \GenStrobeI2C|ALT_INV_ClkCounter\(0),
	datae => \GenStrobeI2C|ALT_INV_ClkCounter\(2),
	dataf => \GenStrobeI2C|ALT_INV_ClkCounter[1]~DUPLICATE_q\,
	combout => \GenStrobeI2C|ClkCounter[2]~3_combout\);

-- Location: FF_X18_Y66_N1
\GenStrobeI2C|ClkCounter[2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \GenStrobeI2C|ClkCounter[2]~3_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \GenStrobeI2C|ClkCounter\(2));

-- Location: LABCELL_X18_Y66_N9
\GenStrobeI2C|ClkCounter[3]~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \GenStrobeI2C|ClkCounter[3]~2_combout\ = ( \GenStrobeI2C|ClkCounter\(3) & ( \GenStrobeI2C|ClkCounter\(2) & ( (!\GenStrobeI2C|ClkCounter\(1)) # (!\GenStrobeI2C|ClkCounter\(0)) ) ) ) # ( !\GenStrobeI2C|ClkCounter\(3) & ( \GenStrobeI2C|ClkCounter\(2) & ( 
-- (\GenStrobeI2C|ClkCounter\(1) & \GenStrobeI2C|ClkCounter\(0)) ) ) ) # ( \GenStrobeI2C|ClkCounter\(3) & ( !\GenStrobeI2C|ClkCounter\(2) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000010101011111111110101010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \GenStrobeI2C|ALT_INV_ClkCounter\(1),
	datad => \GenStrobeI2C|ALT_INV_ClkCounter\(0),
	datae => \GenStrobeI2C|ALT_INV_ClkCounter\(3),
	dataf => \GenStrobeI2C|ALT_INV_ClkCounter\(2),
	combout => \GenStrobeI2C|ClkCounter[3]~2_combout\);

-- Location: FF_X18_Y66_N11
\GenStrobeI2C|ClkCounter[3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \GenStrobeI2C|ClkCounter[3]~2_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \GenStrobeI2C|ClkCounter\(3));

-- Location: LABCELL_X18_Y66_N36
\GenStrobeI2C|ClkCounter[4]~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \GenStrobeI2C|ClkCounter[4]~1_combout\ = ( \GenStrobeI2C|ClkCounter\(4) & ( \GenStrobeI2C|ClkCounter\(2) & ( (!\GenStrobeI2C|ClkCounter\(3)) # ((!\GenStrobeI2C|ClkCounter\(1)) # (!\GenStrobeI2C|ClkCounter[0]~DUPLICATE_q\)) ) ) ) # ( 
-- !\GenStrobeI2C|ClkCounter\(4) & ( \GenStrobeI2C|ClkCounter\(2) & ( (\GenStrobeI2C|ClkCounter\(3) & (\GenStrobeI2C|ClkCounter\(1) & \GenStrobeI2C|ClkCounter[0]~DUPLICATE_q\)) ) ) ) # ( \GenStrobeI2C|ClkCounter\(4) & ( !\GenStrobeI2C|ClkCounter\(2) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000111111111111111100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \GenStrobeI2C|ALT_INV_ClkCounter\(3),
	datac => \GenStrobeI2C|ALT_INV_ClkCounter\(1),
	datad => \GenStrobeI2C|ALT_INV_ClkCounter[0]~DUPLICATE_q\,
	datae => \GenStrobeI2C|ALT_INV_ClkCounter\(4),
	dataf => \GenStrobeI2C|ALT_INV_ClkCounter\(2),
	combout => \GenStrobeI2C|ClkCounter[4]~1_combout\);

-- Location: FF_X18_Y66_N38
\GenStrobeI2C|ClkCounter[4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \GenStrobeI2C|ClkCounter[4]~1_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \GenStrobeI2C|ClkCounter\(4));

-- Location: LABCELL_X18_Y66_N54
\GenStrobeI2C|ClkCounter[5]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \GenStrobeI2C|ClkCounter[5]~0_combout\ = ( \GenStrobeI2C|ClkCounter\(5) & ( \GenStrobeI2C|ClkCounter\(2) & ( (!\GenStrobeI2C|ClkCounter\(4)) # ((!\GenStrobeI2C|ClkCounter[0]~DUPLICATE_q\) # ((!\GenStrobeI2C|ClkCounter[1]~DUPLICATE_q\) # 
-- (!\GenStrobeI2C|ClkCounter\(3)))) ) ) ) # ( !\GenStrobeI2C|ClkCounter\(5) & ( \GenStrobeI2C|ClkCounter\(2) & ( (\GenStrobeI2C|ClkCounter\(4) & (\GenStrobeI2C|ClkCounter[0]~DUPLICATE_q\ & (\GenStrobeI2C|ClkCounter[1]~DUPLICATE_q\ & 
-- \GenStrobeI2C|ClkCounter\(3)))) ) ) ) # ( \GenStrobeI2C|ClkCounter\(5) & ( !\GenStrobeI2C|ClkCounter\(2) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000011111111111111110",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \GenStrobeI2C|ALT_INV_ClkCounter\(4),
	datab => \GenStrobeI2C|ALT_INV_ClkCounter[0]~DUPLICATE_q\,
	datac => \GenStrobeI2C|ALT_INV_ClkCounter[1]~DUPLICATE_q\,
	datad => \GenStrobeI2C|ALT_INV_ClkCounter\(3),
	datae => \GenStrobeI2C|ALT_INV_ClkCounter\(5),
	dataf => \GenStrobeI2C|ALT_INV_ClkCounter\(2),
	combout => \GenStrobeI2C|ClkCounter[5]~0_combout\);

-- Location: FF_X18_Y66_N55
\GenStrobeI2C|ClkCounter[5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \GenStrobeI2C|ClkCounter[5]~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \GenStrobeI2C|ClkCounter\(5));

-- Location: LABCELL_X18_Y66_N12
\GenStrobeI2C|Equal0~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \GenStrobeI2C|Equal0~0_combout\ = ( \GenStrobeI2C|ClkCounter\(5) & ( \GenStrobeI2C|ClkCounter\(2) & ( (\GenStrobeI2C|ClkCounter[1]~DUPLICATE_q\ & (\GenStrobeI2C|ClkCounter[0]~DUPLICATE_q\ & (\GenStrobeI2C|ClkCounter\(4) & \GenStrobeI2C|ClkCounter\(3)))) ) 
-- ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000000000000000000000000001",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \GenStrobeI2C|ALT_INV_ClkCounter[1]~DUPLICATE_q\,
	datab => \GenStrobeI2C|ALT_INV_ClkCounter[0]~DUPLICATE_q\,
	datac => \GenStrobeI2C|ALT_INV_ClkCounter\(4),
	datad => \GenStrobeI2C|ALT_INV_ClkCounter\(3),
	datae => \GenStrobeI2C|ALT_INV_ClkCounter\(5),
	dataf => \GenStrobeI2C|ALT_INV_ClkCounter\(2),
	combout => \GenStrobeI2C|Equal0~0_combout\);

-- Location: FF_X18_Y66_N13
\GenStrobeI2C|oStrobe\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \GenStrobeI2C|Equal0~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \GenStrobeI2C|oStrobe~q\);

-- Location: FF_X19_Y70_N13
\ConfigureCodec|R.FrameState.Idle~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \ConfigureCodec|Selector0~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ConfigureCodec|R.FrameState.Idle~DUPLICATE_q\);

-- Location: MLABCELL_X21_Y70_N0
\ConfigureCodec|Add0~25\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Add0~25_sumout\ = SUM(( \ConfigureCodec|R.AddrCtr\(0) ) + ( VCC ) + ( !VCC ))
-- \ConfigureCodec|Add0~26\ = CARRY(( \ConfigureCodec|R.AddrCtr\(0) ) + ( VCC ) + ( !VCC ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \ConfigureCodec|ALT_INV_R.AddrCtr\(0),
	cin => GND,
	sumout => \ConfigureCodec|Add0~25_sumout\,
	cout => \ConfigureCodec|Add0~26\);

-- Location: FF_X21_Y70_N2
\ConfigureCodec|R.AddrCtr[0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \ConfigureCodec|Add0~25_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \ConfigureCodec|ALT_INV_R.Activity~q\,
	ena => \ConfigureCodec|R.AddrCtr[6]~2_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ConfigureCodec|R.AddrCtr\(0));

-- Location: MLABCELL_X21_Y70_N3
\ConfigureCodec|Add0~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Add0~5_sumout\ = SUM(( \ConfigureCodec|R.AddrCtr\(1) ) + ( GND ) + ( \ConfigureCodec|Add0~26\ ))
-- \ConfigureCodec|Add0~6\ = CARRY(( \ConfigureCodec|R.AddrCtr\(1) ) + ( GND ) + ( \ConfigureCodec|Add0~26\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \ConfigureCodec|ALT_INV_R.AddrCtr\(1),
	cin => \ConfigureCodec|Add0~26\,
	sumout => \ConfigureCodec|Add0~5_sumout\,
	cout => \ConfigureCodec|Add0~6\);

-- Location: FF_X21_Y70_N5
\ConfigureCodec|R.AddrCtr[1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \ConfigureCodec|Add0~5_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \ConfigureCodec|ALT_INV_R.Activity~q\,
	ena => \ConfigureCodec|R.AddrCtr[6]~2_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ConfigureCodec|R.AddrCtr\(1));

-- Location: MLABCELL_X21_Y70_N6
\ConfigureCodec|Add0~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Add0~1_sumout\ = SUM(( \ConfigureCodec|R.AddrCtr\(2) ) + ( GND ) + ( \ConfigureCodec|Add0~6\ ))
-- \ConfigureCodec|Add0~2\ = CARRY(( \ConfigureCodec|R.AddrCtr\(2) ) + ( GND ) + ( \ConfigureCodec|Add0~6\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \ConfigureCodec|ALT_INV_R.AddrCtr\(2),
	cin => \ConfigureCodec|Add0~6\,
	sumout => \ConfigureCodec|Add0~1_sumout\,
	cout => \ConfigureCodec|Add0~2\);

-- Location: MLABCELL_X21_Y70_N9
\ConfigureCodec|Add0~21\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Add0~21_sumout\ = SUM(( \ConfigureCodec|R.AddrCtr\(3) ) + ( GND ) + ( \ConfigureCodec|Add0~2\ ))
-- \ConfigureCodec|Add0~22\ = CARRY(( \ConfigureCodec|R.AddrCtr\(3) ) + ( GND ) + ( \ConfigureCodec|Add0~2\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \ConfigureCodec|ALT_INV_R.AddrCtr\(3),
	cin => \ConfigureCodec|Add0~2\,
	sumout => \ConfigureCodec|Add0~21_sumout\,
	cout => \ConfigureCodec|Add0~22\);

-- Location: FF_X21_Y70_N11
\ConfigureCodec|R.AddrCtr[3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \ConfigureCodec|Add0~21_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \ConfigureCodec|ALT_INV_R.Activity~q\,
	ena => \ConfigureCodec|R.AddrCtr[6]~2_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ConfigureCodec|R.AddrCtr\(3));

-- Location: MLABCELL_X21_Y70_N12
\ConfigureCodec|Add0~17\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Add0~17_sumout\ = SUM(( \ConfigureCodec|R.AddrCtr\(4) ) + ( GND ) + ( \ConfigureCodec|Add0~22\ ))
-- \ConfigureCodec|Add0~18\ = CARRY(( \ConfigureCodec|R.AddrCtr\(4) ) + ( GND ) + ( \ConfigureCodec|Add0~22\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \ConfigureCodec|ALT_INV_R.AddrCtr\(4),
	cin => \ConfigureCodec|Add0~22\,
	sumout => \ConfigureCodec|Add0~17_sumout\,
	cout => \ConfigureCodec|Add0~18\);

-- Location: FF_X21_Y70_N14
\ConfigureCodec|R.AddrCtr[4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \ConfigureCodec|Add0~17_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \ConfigureCodec|ALT_INV_R.Activity~q\,
	ena => \ConfigureCodec|R.AddrCtr[6]~2_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ConfigureCodec|R.AddrCtr\(4));

-- Location: MLABCELL_X21_Y70_N15
\ConfigureCodec|Add0~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Add0~13_sumout\ = SUM(( \ConfigureCodec|R.AddrCtr\(5) ) + ( GND ) + ( \ConfigureCodec|Add0~18\ ))
-- \ConfigureCodec|Add0~14\ = CARRY(( \ConfigureCodec|R.AddrCtr\(5) ) + ( GND ) + ( \ConfigureCodec|Add0~18\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \ConfigureCodec|ALT_INV_R.AddrCtr\(5),
	cin => \ConfigureCodec|Add0~18\,
	sumout => \ConfigureCodec|Add0~13_sumout\,
	cout => \ConfigureCodec|Add0~14\);

-- Location: FF_X21_Y70_N17
\ConfigureCodec|R.AddrCtr[5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \ConfigureCodec|Add0~13_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \ConfigureCodec|ALT_INV_R.Activity~q\,
	ena => \ConfigureCodec|R.AddrCtr[6]~2_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ConfigureCodec|R.AddrCtr\(5));

-- Location: MLABCELL_X21_Y70_N18
\ConfigureCodec|Add0~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Add0~9_sumout\ = SUM(( \ConfigureCodec|R.AddrCtr\(6) ) + ( GND ) + ( \ConfigureCodec|Add0~14\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \ConfigureCodec|ALT_INV_R.AddrCtr\(6),
	cin => \ConfigureCodec|Add0~14\,
	sumout => \ConfigureCodec|Add0~9_sumout\);

-- Location: FF_X21_Y70_N20
\ConfigureCodec|R.AddrCtr[6]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \ConfigureCodec|Add0~9_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \ConfigureCodec|ALT_INV_R.Activity~q\,
	ena => \ConfigureCodec|R.AddrCtr[6]~2_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ConfigureCodec|R.AddrCtr\(6));

-- Location: MLABCELL_X21_Y70_N48
\ConfigureCodec|Equal0~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Equal0~1_combout\ = ( !\ConfigureCodec|R.AddrCtr\(5) & ( (\ConfigureCodec|R.AddrCtr\(0) & (\ConfigureCodec|R.AddrCtr\(3) & (!\ConfigureCodec|R.AddrCtr\(6) & !\ConfigureCodec|R.AddrCtr\(4)))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000000000000000100000000000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ConfigureCodec|ALT_INV_R.AddrCtr\(0),
	datab => \ConfigureCodec|ALT_INV_R.AddrCtr\(3),
	datac => \ConfigureCodec|ALT_INV_R.AddrCtr\(6),
	datad => \ConfigureCodec|ALT_INV_R.AddrCtr\(4),
	dataf => \ConfigureCodec|ALT_INV_R.AddrCtr\(5),
	combout => \ConfigureCodec|Equal0~1_combout\);

-- Location: LABCELL_X19_Y70_N21
\ConfigureCodec|Selector1~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Selector1~1_combout\ = ( \ConfigureCodec|R.Activity~q\ & ( (!\GenStrobeI2C|oStrobe~q\ & ((\ConfigureCodec|R.FrameState.Start~q\))) # (\GenStrobeI2C|oStrobe~q\ & (!\ConfigureCodec|R.FrameState.Idle~q\)) ) ) # ( 
-- !\ConfigureCodec|R.Activity~q\ & ( (!\GenStrobeI2C|oStrobe~q\ & \ConfigureCodec|R.FrameState.Start~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000010101010000000001010101001010000111110100101000011111010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \GenStrobeI2C|ALT_INV_oStrobe~q\,
	datac => \ConfigureCodec|ALT_INV_R.FrameState.Idle~q\,
	datad => \ConfigureCodec|ALT_INV_R.FrameState.Start~q\,
	dataf => \ConfigureCodec|ALT_INV_R.Activity~q\,
	combout => \ConfigureCodec|Selector1~1_combout\);

-- Location: FF_X19_Y70_N22
\ConfigureCodec|R.FrameState.Start\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \ConfigureCodec|Selector1~1_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ConfigureCodec|R.FrameState.Start~q\);

-- Location: LABCELL_X17_Y70_N51
\ConfigureCodec|Selector1~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Selector1~0_combout\ = (\ConfigureCodec|R.FrameState.Start~q\ & !\GenStrobeI2C|oStrobe~q\)

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011000000110000001100000011000000110000001100000011000000110000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ConfigureCodec|ALT_INV_R.FrameState.Start~q\,
	datac => \GenStrobeI2C|ALT_INV_oStrobe~q\,
	combout => \ConfigureCodec|Selector1~0_combout\);

-- Location: LABCELL_X17_Y70_N15
\ConfigureCodec|NextStateAndOutput:vSclkFalling~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|NextStateAndOutput:vSclkFalling~0_combout\ = ( !\ConfigureCodec|R.Sclk~q\ & ( \GenStrobeI2C|oStrobe~q\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111000000000000000000001111000011110000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \GenStrobeI2C|ALT_INV_oStrobe~q\,
	datae => \ConfigureCodec|ALT_INV_R.Sclk~q\,
	combout => \ConfigureCodec|NextStateAndOutput:vSclkFalling~0_combout\);

-- Location: FF_X18_Y70_N49
\ConfigureCodec|R.BitCtr[3]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \ConfigureCodec|Selector10~2_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ConfigureCodec|R.BitCtr[3]~DUPLICATE_q\);

-- Location: LABCELL_X19_Y70_N27
\ConfigureCodec|Selector2~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Selector2~0_combout\ = ( \ConfigureCodec|R.FrameState.Start~q\ & ( ((!\ConfigureCodec|NextR~8_combout\ & \ConfigureCodec|R.FrameState.Address~q\)) # (\GenStrobeI2C|oStrobe~q\) ) ) # ( !\ConfigureCodec|R.FrameState.Start~q\ & ( 
-- (!\ConfigureCodec|NextR~8_combout\ & \ConfigureCodec|R.FrameState.Address~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011110000000000001111000001010101111101010101010111110101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \GenStrobeI2C|ALT_INV_oStrobe~q\,
	datac => \ConfigureCodec|ALT_INV_NextR~8_combout\,
	datad => \ConfigureCodec|ALT_INV_R.FrameState.Address~q\,
	dataf => \ConfigureCodec|ALT_INV_R.FrameState.Start~q\,
	combout => \ConfigureCodec|Selector2~0_combout\);

-- Location: FF_X19_Y70_N28
\ConfigureCodec|R.FrameState.Address\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \ConfigureCodec|Selector2~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ConfigureCodec|R.FrameState.Address~q\);

-- Location: LABCELL_X19_Y70_N36
\ConfigureCodec|Selector3~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Selector3~0_combout\ = ( \ConfigureCodec|R.FrameState.Address~q\ & ( ((!\ConfigureCodec|NextStateAndOutput:vSclkFalling~0_combout\ & \ConfigureCodec|R.FrameState.RWBit~q\)) # (\ConfigureCodec|NextR~8_combout\) ) ) # ( 
-- !\ConfigureCodec|R.FrameState.Address~q\ & ( (!\ConfigureCodec|NextStateAndOutput:vSclkFalling~0_combout\ & \ConfigureCodec|R.FrameState.RWBit~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011110000000000001111000000110011111100110011001111110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ConfigureCodec|ALT_INV_NextR~8_combout\,
	datac => \ConfigureCodec|ALT_INV_NextStateAndOutput:vSclkFalling~0_combout\,
	datad => \ConfigureCodec|ALT_INV_R.FrameState.RWBit~q\,
	dataf => \ConfigureCodec|ALT_INV_R.FrameState.Address~q\,
	combout => \ConfigureCodec|Selector3~0_combout\);

-- Location: FF_X19_Y70_N37
\ConfigureCodec|R.FrameState.RWBit\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \ConfigureCodec|Selector3~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ConfigureCodec|R.FrameState.RWBit~q\);

-- Location: FF_X19_Y70_N41
\ConfigureCodec|R.FrameState.Ack1\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \ConfigureCodec|R.FrameState.Ack1~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ConfigureCodec|R.FrameState.Ack1~q\);

-- Location: LABCELL_X19_Y70_N39
\ConfigureCodec|R.FrameState.Ack1~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|R.FrameState.Ack1~0_combout\ = ( \ConfigureCodec|R.Sclk~q\ & ( \ConfigureCodec|R.FrameState.Ack1~q\ ) ) # ( !\ConfigureCodec|R.Sclk~q\ & ( (!\GenStrobeI2C|oStrobe~q\ & ((\ConfigureCodec|R.FrameState.Ack1~q\))) # (\GenStrobeI2C|oStrobe~q\ & 
-- (\ConfigureCodec|R.FrameState.RWBit~q\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010110101111000001011010111100000000111111110000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \GenStrobeI2C|ALT_INV_oStrobe~q\,
	datac => \ConfigureCodec|ALT_INV_R.FrameState.RWBit~q\,
	datad => \ConfigureCodec|ALT_INV_R.FrameState.Ack1~q\,
	dataf => \ConfigureCodec|ALT_INV_R.Sclk~q\,
	combout => \ConfigureCodec|R.FrameState.Ack1~0_combout\);

-- Location: FF_X19_Y70_N40
\ConfigureCodec|R.FrameState.Ack1~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \ConfigureCodec|R.FrameState.Ack1~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ConfigureCodec|R.FrameState.Ack1~DUPLICATE_q\);

-- Location: LABCELL_X19_Y70_N45
\ConfigureCodec|Selector8~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Selector8~0_combout\ = ( \ConfigureCodec|R.FrameState.Data2~DUPLICATE_q\ & ( ((!\ConfigureCodec|NextStateAndOutput:vSclkFalling~0_combout\ & \ConfigureCodec|R.FrameState.Ack3~q\)) # (\ConfigureCodec|NextR~8_combout\) ) ) # ( 
-- !\ConfigureCodec|R.FrameState.Data2~DUPLICATE_q\ & ( (!\ConfigureCodec|NextStateAndOutput:vSclkFalling~0_combout\ & \ConfigureCodec|R.FrameState.Ack3~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011001100000000001100110000001111110011110000111111001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ConfigureCodec|ALT_INV_NextStateAndOutput:vSclkFalling~0_combout\,
	datac => \ConfigureCodec|ALT_INV_NextR~8_combout\,
	datad => \ConfigureCodec|ALT_INV_R.FrameState.Ack3~q\,
	dataf => \ConfigureCodec|ALT_INV_R.FrameState.Data2~DUPLICATE_q\,
	combout => \ConfigureCodec|Selector8~0_combout\);

-- Location: FF_X19_Y70_N46
\ConfigureCodec|R.FrameState.Ack3\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \ConfigureCodec|Selector8~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ConfigureCodec|R.FrameState.Ack3~q\);

-- Location: LABCELL_X19_Y70_N33
\ConfigureCodec|Selector13~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Selector13~0_combout\ = ( !\ConfigureCodec|R.FrameState.Ack1~q\ & ( (!\ConfigureCodec|R.FrameState.Ack2~q\ & !\ConfigureCodec|R.FrameState.Ack3~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1010000010100000101000001010000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ConfigureCodec|ALT_INV_R.FrameState.Ack2~q\,
	datac => \ConfigureCodec|ALT_INV_R.FrameState.Ack3~q\,
	dataf => \ConfigureCodec|ALT_INV_R.FrameState.Ack1~q\,
	combout => \ConfigureCodec|Selector13~0_combout\);

-- Location: IOIBUF_X12_Y81_N1
\ioI2cSdin~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ioI2cSdin,
	o => \ioI2cSdin~input_o\);

-- Location: LABCELL_X19_Y70_N48
\ConfigureCodec|Selector16~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Selector16~1_combout\ = ( \ConfigureCodec|R.AckError~q\ & ( \ConfigureCodec|R.Sclk~q\ & ( (!\GenStrobeI2C|oStrobe~q\) # ((!\ConfigureCodec|R.AddrCtr[6]~0_combout\) # ((!\ConfigureCodec|Selector13~0_combout\ & \ioI2cSdin~input_o\))) ) ) ) # 
-- ( !\ConfigureCodec|R.AckError~q\ & ( \ConfigureCodec|R.Sclk~q\ & ( (\GenStrobeI2C|oStrobe~q\ & (!\ConfigureCodec|Selector13~0_combout\ & \ioI2cSdin~input_o\)) ) ) ) # ( \ConfigureCodec|R.AckError~q\ & ( !\ConfigureCodec|R.Sclk~q\ & ( 
-- (!\GenStrobeI2C|oStrobe~q\) # (!\ConfigureCodec|R.AddrCtr[6]~0_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111011101110111000000000010100001110111011111110",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \GenStrobeI2C|ALT_INV_oStrobe~q\,
	datab => \ConfigureCodec|ALT_INV_R.AddrCtr[6]~0_combout\,
	datac => \ConfigureCodec|ALT_INV_Selector13~0_combout\,
	datad => \ALT_INV_ioI2cSdin~input_o\,
	datae => \ConfigureCodec|ALT_INV_R.AckError~q\,
	dataf => \ConfigureCodec|ALT_INV_R.Sclk~q\,
	combout => \ConfigureCodec|Selector16~1_combout\);

-- Location: FF_X19_Y70_N50
\ConfigureCodec|R.AckError\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \ConfigureCodec|Selector16~1_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ConfigureCodec|R.AckError~q\);

-- Location: LABCELL_X17_Y70_N48
\ConfigureCodec|Selector5~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Selector5~0_combout\ = (!\ConfigureCodec|R.AckError~q\ & \ConfigureCodec|R.FrameState.Ack1~DUPLICATE_q\)

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000101000001010000010100000101000001010000010100000101000001010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ConfigureCodec|ALT_INV_R.AckError~q\,
	datac => \ConfigureCodec|ALT_INV_R.FrameState.Ack1~DUPLICATE_q\,
	combout => \ConfigureCodec|Selector5~0_combout\);

-- Location: FF_X18_Y70_N37
\ConfigureCodec|R.FrameState.Data1\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \ConfigureCodec|Selector5~1_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ConfigureCodec|R.FrameState.Data1~q\);

-- Location: LABCELL_X18_Y70_N36
\ConfigureCodec|Selector5~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Selector5~1_combout\ = ( \ConfigureCodec|NextR~9_combout\ & ( (!\ConfigureCodec|NextStateAndOutput:vSclkFalling~0_combout\ & (((\ConfigureCodec|R.FrameState.Data1~q\)))) # (\ConfigureCodec|NextStateAndOutput:vSclkFalling~0_combout\ & 
-- (((!\ConfigureCodec|R.BitCtr\(3) & \ConfigureCodec|R.FrameState.Data1~q\)) # (\ConfigureCodec|Selector5~0_combout\))) ) ) # ( !\ConfigureCodec|NextR~9_combout\ & ( ((\ConfigureCodec|NextStateAndOutput:vSclkFalling~0_combout\ & 
-- \ConfigureCodec|Selector5~0_combout\)) # (\ConfigureCodec|R.FrameState.Data1~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001111111111000000111111111100000011111011110000001111101111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ConfigureCodec|ALT_INV_R.BitCtr\(3),
	datab => \ConfigureCodec|ALT_INV_NextStateAndOutput:vSclkFalling~0_combout\,
	datac => \ConfigureCodec|ALT_INV_Selector5~0_combout\,
	datad => \ConfigureCodec|ALT_INV_R.FrameState.Data1~q\,
	dataf => \ConfigureCodec|ALT_INV_NextR~9_combout\,
	combout => \ConfigureCodec|Selector5~1_combout\);

-- Location: FF_X18_Y70_N38
\ConfigureCodec|R.FrameState.Data1~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \ConfigureCodec|Selector5~1_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ConfigureCodec|R.FrameState.Data1~DUPLICATE_q\);

-- Location: LABCELL_X17_Y70_N54
\ConfigureCodec|Selector13~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Selector13~2_combout\ = ( \ConfigureCodec|R.BitCtr\(0) & ( \GenStrobeI2C|oStrobe~q\ & ( (!\ConfigureCodec|R.Sclk~q\ & (\ConfigureCodec|R.FrameState.Ack1~DUPLICATE_q\ & ((!\ConfigureCodec|R.AckError~q\)))) # (\ConfigureCodec|R.Sclk~q\ & 
-- (((\ConfigureCodec|R.FrameState.Data1~DUPLICATE_q\)))) ) ) ) # ( !\ConfigureCodec|R.BitCtr\(0) & ( \GenStrobeI2C|oStrobe~q\ & ( (!\ConfigureCodec|R.Sclk~q\ & (((\ConfigureCodec|R.FrameState.Ack1~DUPLICATE_q\ & !\ConfigureCodec|R.AckError~q\)) # 
-- (\ConfigureCodec|R.FrameState.Data1~DUPLICATE_q\))) ) ) ) # ( \ConfigureCodec|R.BitCtr\(0) & ( !\GenStrobeI2C|oStrobe~q\ & ( \ConfigureCodec|R.FrameState.Data1~DUPLICATE_q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000001100110011001101110011000000000101000000110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ConfigureCodec|ALT_INV_R.FrameState.Ack1~DUPLICATE_q\,
	datab => \ConfigureCodec|ALT_INV_R.FrameState.Data1~DUPLICATE_q\,
	datac => \ConfigureCodec|ALT_INV_R.AckError~q\,
	datad => \ConfigureCodec|ALT_INV_R.Sclk~q\,
	datae => \ConfigureCodec|ALT_INV_R.BitCtr\(0),
	dataf => \GenStrobeI2C|ALT_INV_oStrobe~q\,
	combout => \ConfigureCodec|Selector13~2_combout\);

-- Location: LABCELL_X19_Y70_N6
\ConfigureCodec|Selector13~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Selector13~1_combout\ = ( !\ConfigureCodec|R.FrameState.RWBit~q\ & ( \ConfigureCodec|R.FrameState.Idle~q\ & ( (!\ConfigureCodec|R.FrameState.Stop~q\ & (!\ConfigureCodec|R.FrameState.Ack1~q\ & (!\ConfigureCodec|R.FrameState.Ack2~q\ & 
-- !\ConfigureCodec|R.FrameState.Ack3~q\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000010000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ConfigureCodec|ALT_INV_R.FrameState.Stop~q\,
	datab => \ConfigureCodec|ALT_INV_R.FrameState.Ack1~q\,
	datac => \ConfigureCodec|ALT_INV_R.FrameState.Ack2~q\,
	datad => \ConfigureCodec|ALT_INV_R.FrameState.Ack3~q\,
	datae => \ConfigureCodec|ALT_INV_R.FrameState.RWBit~q\,
	dataf => \ConfigureCodec|ALT_INV_R.FrameState.Idle~q\,
	combout => \ConfigureCodec|Selector13~1_combout\);

-- Location: LABCELL_X17_Y70_N24
\ConfigureCodec|NextR~10\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|NextR~10_combout\ = ( \ConfigureCodec|R.BitCtr\(0) & ( \GenStrobeI2C|oStrobe~q\ & ( !\ConfigureCodec|R.Sclk~q\ ) ) ) # ( !\ConfigureCodec|R.BitCtr\(0) & ( \GenStrobeI2C|oStrobe~q\ & ( (!\ConfigureCodec|R.Sclk~q\ & 
-- (((\ConfigureCodec|R.BitCtr\(1)) # (\ConfigureCodec|R.BitCtr\(2))) # (\ConfigureCodec|R.BitCtr[3]~DUPLICATE_q\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000001001100110011001100110011001100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ConfigureCodec|ALT_INV_R.BitCtr[3]~DUPLICATE_q\,
	datab => \ConfigureCodec|ALT_INV_R.Sclk~q\,
	datac => \ConfigureCodec|ALT_INV_R.BitCtr\(2),
	datad => \ConfigureCodec|ALT_INV_R.BitCtr\(1),
	datae => \ConfigureCodec|ALT_INV_R.BitCtr\(0),
	dataf => \GenStrobeI2C|ALT_INV_oStrobe~q\,
	combout => \ConfigureCodec|NextR~10_combout\);

-- Location: LABCELL_X17_Y70_N0
\ConfigureCodec|Selector13~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Selector13~3_combout\ = ( \ConfigureCodec|R.BitCtr\(0) & ( \ConfigureCodec|NextR~10_combout\ & ( ((!\ConfigureCodec|Selector13~1_combout\) # (\ConfigureCodec|Selector13~2_combout\)) # (\ConfigureCodec|Selector1~0_combout\) ) ) ) # ( 
-- !\ConfigureCodec|R.BitCtr\(0) & ( \ConfigureCodec|NextR~10_combout\ & ( (!\ConfigureCodec|Selector10~0_combout\) # (\ConfigureCodec|Selector13~2_combout\) ) ) ) # ( \ConfigureCodec|R.BitCtr\(0) & ( !\ConfigureCodec|NextR~10_combout\ & ( 
-- (!\ConfigureCodec|Selector10~0_combout\) # (((!\ConfigureCodec|Selector13~1_combout\) # (\ConfigureCodec|Selector13~2_combout\)) # (\ConfigureCodec|Selector1~0_combout\)) ) ) ) # ( !\ConfigureCodec|R.BitCtr\(0) & ( !\ConfigureCodec|NextR~10_combout\ & ( 
-- \ConfigureCodec|Selector13~2_combout\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111111111111011111110101111101011111111111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ConfigureCodec|ALT_INV_Selector10~0_combout\,
	datab => \ConfigureCodec|ALT_INV_Selector1~0_combout\,
	datac => \ConfigureCodec|ALT_INV_Selector13~2_combout\,
	datad => \ConfigureCodec|ALT_INV_Selector13~1_combout\,
	datae => \ConfigureCodec|ALT_INV_R.BitCtr\(0),
	dataf => \ConfigureCodec|ALT_INV_NextR~10_combout\,
	combout => \ConfigureCodec|Selector13~3_combout\);

-- Location: FF_X17_Y70_N2
\ConfigureCodec|R.BitCtr[0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \ConfigureCodec|Selector13~3_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ConfigureCodec|R.BitCtr\(0));

-- Location: LABCELL_X17_Y70_N33
\ConfigureCodec|Mux8~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Mux8~0_combout\ = (!\ConfigureCodec|R.BitCtr\(0) & !\ConfigureCodec|R.BitCtr\(1))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1000100010001000100010001000100010001000100010001000100010001000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ConfigureCodec|ALT_INV_R.BitCtr\(0),
	datab => \ConfigureCodec|ALT_INV_R.BitCtr\(1),
	combout => \ConfigureCodec|Mux8~0_combout\);

-- Location: LABCELL_X17_Y70_N42
\ConfigureCodec|Selector11~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Selector11~2_combout\ = ( \ConfigureCodec|R.BitCtr\(2) & ( \ConfigureCodec|Selector10~0_combout\ & ( (\ConfigureCodec|R.FrameState.Start~q\ & \GenStrobeI2C|oStrobe~q\) ) ) ) # ( !\ConfigureCodec|R.BitCtr\(2) & ( 
-- \ConfigureCodec|Selector10~0_combout\ & ( (\ConfigureCodec|R.FrameState.Start~q\ & \GenStrobeI2C|oStrobe~q\) ) ) ) # ( \ConfigureCodec|R.BitCtr\(2) & ( !\ConfigureCodec|Selector10~0_combout\ & ( (!\ConfigureCodec|Mux8~0_combout\) # 
-- ((!\ConfigureCodec|NextR~10_combout\) # ((\ConfigureCodec|R.FrameState.Start~q\ & \GenStrobeI2C|oStrobe~q\))) ) ) ) # ( !\ConfigureCodec|R.BitCtr\(2) & ( !\ConfigureCodec|Selector10~0_combout\ & ( (!\ConfigureCodec|Mux8~0_combout\ & 
-- (\ConfigureCodec|R.FrameState.Start~q\ & ((\GenStrobeI2C|oStrobe~q\)))) # (\ConfigureCodec|Mux8~0_combout\ & (((\ConfigureCodec|R.FrameState.Start~q\ & \GenStrobeI2C|oStrobe~q\)) # (\ConfigureCodec|NextR~10_combout\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100110111111110101111101100000000001100110000000000110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ConfigureCodec|ALT_INV_Mux8~0_combout\,
	datab => \ConfigureCodec|ALT_INV_R.FrameState.Start~q\,
	datac => \ConfigureCodec|ALT_INV_NextR~10_combout\,
	datad => \GenStrobeI2C|ALT_INV_oStrobe~q\,
	datae => \ConfigureCodec|ALT_INV_R.BitCtr\(2),
	dataf => \ConfigureCodec|ALT_INV_Selector10~0_combout\,
	combout => \ConfigureCodec|Selector11~2_combout\);

-- Location: FF_X17_Y70_N1
\ConfigureCodec|R.BitCtr[0]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \ConfigureCodec|Selector13~3_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ConfigureCodec|R.BitCtr[0]~DUPLICATE_q\);

-- Location: LABCELL_X18_Y70_N45
\ConfigureCodec|Selector11~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Selector11~1_combout\ = ( \ConfigureCodec|R.BitCtr\(1) & ( (\ConfigureCodec|R.FrameState.Data1~q\ & \ConfigureCodec|R.BitCtr\(2)) ) ) # ( !\ConfigureCodec|R.BitCtr\(1) & ( (\ConfigureCodec|R.FrameState.Data1~q\ & 
-- (!\ConfigureCodec|R.BitCtr\(2) $ (\ConfigureCodec|R.BitCtr[0]~DUPLICATE_q\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101000000000101010100000000010100000101000001010000010100000101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ConfigureCodec|ALT_INV_R.FrameState.Data1~q\,
	datac => \ConfigureCodec|ALT_INV_R.BitCtr\(2),
	datad => \ConfigureCodec|ALT_INV_R.BitCtr[0]~DUPLICATE_q\,
	dataf => \ConfigureCodec|ALT_INV_R.BitCtr\(1),
	combout => \ConfigureCodec|Selector11~1_combout\);

-- Location: LABCELL_X18_Y70_N27
\ConfigureCodec|Selector11~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Selector11~0_combout\ = ( \ConfigureCodec|R.FrameState.Data1~q\ & ( (\ConfigureCodec|Selector13~1_combout\ & (\ConfigureCodec|NextStateAndOutput:vSclkFalling~0_combout\ & !\ConfigureCodec|R.FrameState.Start~q\)) ) ) # ( 
-- !\ConfigureCodec|R.FrameState.Data1~q\ & ( (\ConfigureCodec|Selector13~1_combout\ & !\ConfigureCodec|R.FrameState.Start~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010100000000010101010000000000000101000000000000010100000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ConfigureCodec|ALT_INV_Selector13~1_combout\,
	datac => \ConfigureCodec|ALT_INV_NextStateAndOutput:vSclkFalling~0_combout\,
	datad => \ConfigureCodec|ALT_INV_R.FrameState.Start~q\,
	dataf => \ConfigureCodec|ALT_INV_R.FrameState.Data1~q\,
	combout => \ConfigureCodec|Selector11~0_combout\);

-- Location: LABCELL_X18_Y70_N54
\ConfigureCodec|Selector11~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Selector11~3_combout\ = ( \ConfigureCodec|R.BitCtr\(2) & ( \ConfigureCodec|Selector11~0_combout\ & ( ((\ConfigureCodec|NextStateAndOutput:vSclkFalling~0_combout\ & ((\ConfigureCodec|Selector11~1_combout\) # 
-- (\ConfigureCodec|Selector5~0_combout\)))) # (\ConfigureCodec|Selector11~2_combout\) ) ) ) # ( !\ConfigureCodec|R.BitCtr\(2) & ( \ConfigureCodec|Selector11~0_combout\ & ( ((\ConfigureCodec|NextStateAndOutput:vSclkFalling~0_combout\ & 
-- ((\ConfigureCodec|Selector11~1_combout\) # (\ConfigureCodec|Selector5~0_combout\)))) # (\ConfigureCodec|Selector11~2_combout\) ) ) ) # ( \ConfigureCodec|R.BitCtr\(2) & ( !\ConfigureCodec|Selector11~0_combout\ ) ) # ( !\ConfigureCodec|R.BitCtr\(2) & ( 
-- !\ConfigureCodec|Selector11~0_combout\ & ( ((\ConfigureCodec|NextStateAndOutput:vSclkFalling~0_combout\ & ((\ConfigureCodec|Selector11~1_combout\) # (\ConfigureCodec|Selector5~0_combout\)))) # (\ConfigureCodec|Selector11~2_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101011101110111111111111111111101010111011101110101011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ConfigureCodec|ALT_INV_Selector11~2_combout\,
	datab => \ConfigureCodec|ALT_INV_NextStateAndOutput:vSclkFalling~0_combout\,
	datac => \ConfigureCodec|ALT_INV_Selector5~0_combout\,
	datad => \ConfigureCodec|ALT_INV_Selector11~1_combout\,
	datae => \ConfigureCodec|ALT_INV_R.BitCtr\(2),
	dataf => \ConfigureCodec|ALT_INV_Selector11~0_combout\,
	combout => \ConfigureCodec|Selector11~3_combout\);

-- Location: FF_X18_Y70_N55
\ConfigureCodec|R.BitCtr[2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \ConfigureCodec|Selector11~3_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ConfigureCodec|R.BitCtr\(2));

-- Location: LABCELL_X17_Y70_N6
\ConfigureCodec|NextR~8\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|NextR~8_combout\ = ( !\ConfigureCodec|R.BitCtr\(0) & ( \GenStrobeI2C|oStrobe~q\ & ( (!\ConfigureCodec|R.BitCtr[3]~DUPLICATE_q\ & (!\ConfigureCodec|R.Sclk~q\ & (!\ConfigureCodec|R.BitCtr\(2) & !\ConfigureCodec|R.BitCtr\(1)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000010000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ConfigureCodec|ALT_INV_R.BitCtr[3]~DUPLICATE_q\,
	datab => \ConfigureCodec|ALT_INV_R.Sclk~q\,
	datac => \ConfigureCodec|ALT_INV_R.BitCtr\(2),
	datad => \ConfigureCodec|ALT_INV_R.BitCtr\(1),
	datae => \ConfigureCodec|ALT_INV_R.BitCtr\(0),
	dataf => \GenStrobeI2C|ALT_INV_oStrobe~q\,
	combout => \ConfigureCodec|NextR~8_combout\);

-- Location: FF_X19_Y70_N32
\ConfigureCodec|R.FrameState.Data2\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \ConfigureCodec|Selector7~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ConfigureCodec|R.FrameState.Data2~q\);

-- Location: LABCELL_X19_Y70_N30
\ConfigureCodec|Selector7~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Selector7~0_combout\ = ( \ConfigureCodec|R.AckError~q\ & ( (!\ConfigureCodec|NextR~8_combout\ & \ConfigureCodec|R.FrameState.Data2~q\) ) ) # ( !\ConfigureCodec|R.AckError~q\ & ( (!\ConfigureCodec|R.FrameState.Ack2~q\ & 
-- (((!\ConfigureCodec|NextR~8_combout\ & \ConfigureCodec|R.FrameState.Data2~q\)))) # (\ConfigureCodec|R.FrameState.Ack2~q\ & (((!\ConfigureCodec|NextR~8_combout\ & \ConfigureCodec|R.FrameState.Data2~q\)) # 
-- (\ConfigureCodec|NextStateAndOutput:vSclkFalling~0_combout\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000111110001000100011111000100000000111100000000000011110000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ConfigureCodec|ALT_INV_R.FrameState.Ack2~q\,
	datab => \ConfigureCodec|ALT_INV_NextStateAndOutput:vSclkFalling~0_combout\,
	datac => \ConfigureCodec|ALT_INV_NextR~8_combout\,
	datad => \ConfigureCodec|ALT_INV_R.FrameState.Data2~q\,
	dataf => \ConfigureCodec|ALT_INV_R.AckError~q\,
	combout => \ConfigureCodec|Selector7~0_combout\);

-- Location: FF_X19_Y70_N31
\ConfigureCodec|R.FrameState.Data2~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \ConfigureCodec|Selector7~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ConfigureCodec|R.FrameState.Data2~DUPLICATE_q\);

-- Location: LABCELL_X19_Y70_N42
\ConfigureCodec|Selector10~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Selector10~0_combout\ = ( !\ConfigureCodec|R.FrameState.Address~q\ & ( !\ConfigureCodec|R.FrameState.Data2~DUPLICATE_q\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1010101010101010101010101010101000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ConfigureCodec|ALT_INV_R.FrameState.Data2~DUPLICATE_q\,
	dataf => \ConfigureCodec|ALT_INV_R.FrameState.Address~q\,
	combout => \ConfigureCodec|Selector10~0_combout\);

-- Location: LABCELL_X17_Y70_N36
\ConfigureCodec|Selector12~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Selector12~1_combout\ = ( \ConfigureCodec|R.FrameState.Start~q\ & ( \ConfigureCodec|NextR~10_combout\ & ( ((!\ConfigureCodec|Selector10~0_combout\ & (!\ConfigureCodec|R.BitCtr\(1) $ (\ConfigureCodec|R.BitCtr\(0))))) # 
-- (\GenStrobeI2C|oStrobe~q\) ) ) ) # ( !\ConfigureCodec|R.FrameState.Start~q\ & ( \ConfigureCodec|NextR~10_combout\ & ( (!\ConfigureCodec|Selector10~0_combout\ & (!\ConfigureCodec|R.BitCtr\(1) $ (\ConfigureCodec|R.BitCtr\(0)))) ) ) ) # ( 
-- \ConfigureCodec|R.FrameState.Start~q\ & ( !\ConfigureCodec|NextR~10_combout\ & ( ((!\ConfigureCodec|Selector10~0_combout\ & \ConfigureCodec|R.BitCtr\(1))) # (\GenStrobeI2C|oStrobe~q\) ) ) ) # ( !\ConfigureCodec|R.FrameState.Start~q\ & ( 
-- !\ConfigureCodec|NextR~10_combout\ & ( (!\ConfigureCodec|Selector10~0_combout\ & \ConfigureCodec|R.BitCtr\(1)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0010001000100010001000101111111110000010100000101000001011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ConfigureCodec|ALT_INV_Selector10~0_combout\,
	datab => \ConfigureCodec|ALT_INV_R.BitCtr\(1),
	datac => \ConfigureCodec|ALT_INV_R.BitCtr\(0),
	datad => \GenStrobeI2C|ALT_INV_oStrobe~q\,
	datae => \ConfigureCodec|ALT_INV_R.FrameState.Start~q\,
	dataf => \ConfigureCodec|ALT_INV_NextR~10_combout\,
	combout => \ConfigureCodec|Selector12~1_combout\);

-- Location: LABCELL_X17_Y70_N30
\ConfigureCodec|Selector12~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Selector12~0_combout\ = ( \ConfigureCodec|R.FrameState.Ack1~DUPLICATE_q\ & ( (!\ConfigureCodec|R.AckError~q\) # ((\ConfigureCodec|R.FrameState.Data1~DUPLICATE_q\ & (!\ConfigureCodec|R.BitCtr\(0) $ (\ConfigureCodec|R.BitCtr\(1))))) ) ) # ( 
-- !\ConfigureCodec|R.FrameState.Ack1~DUPLICATE_q\ & ( (\ConfigureCodec|R.FrameState.Data1~DUPLICATE_q\ & (!\ConfigureCodec|R.BitCtr\(0) $ (\ConfigureCodec|R.BitCtr\(1)))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000010011001000000001001100111110000111110011111000011111001",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ConfigureCodec|ALT_INV_R.BitCtr\(0),
	datab => \ConfigureCodec|ALT_INV_R.BitCtr\(1),
	datac => \ConfigureCodec|ALT_INV_R.AckError~q\,
	datad => \ConfigureCodec|ALT_INV_R.FrameState.Data1~DUPLICATE_q\,
	dataf => \ConfigureCodec|ALT_INV_R.FrameState.Ack1~DUPLICATE_q\,
	combout => \ConfigureCodec|Selector12~0_combout\);

-- Location: LABCELL_X17_Y70_N18
\ConfigureCodec|Selector12~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Selector12~2_combout\ = ( \ConfigureCodec|R.BitCtr\(1) & ( \ConfigureCodec|Selector12~0_combout\ & ( ((!\ConfigureCodec|Selector11~0_combout\) # (\ConfigureCodec|NextStateAndOutput:vSclkFalling~0_combout\)) # 
-- (\ConfigureCodec|Selector12~1_combout\) ) ) ) # ( !\ConfigureCodec|R.BitCtr\(1) & ( \ConfigureCodec|Selector12~0_combout\ & ( (\ConfigureCodec|NextStateAndOutput:vSclkFalling~0_combout\) # (\ConfigureCodec|Selector12~1_combout\) ) ) ) # ( 
-- \ConfigureCodec|R.BitCtr\(1) & ( !\ConfigureCodec|Selector12~0_combout\ & ( (!\ConfigureCodec|Selector11~0_combout\) # (\ConfigureCodec|Selector12~1_combout\) ) ) ) # ( !\ConfigureCodec|R.BitCtr\(1) & ( !\ConfigureCodec|Selector12~0_combout\ & ( 
-- \ConfigureCodec|Selector12~1_combout\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010101010101111101011111010101110111011101111111011111110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ConfigureCodec|ALT_INV_Selector12~1_combout\,
	datab => \ConfigureCodec|ALT_INV_NextStateAndOutput:vSclkFalling~0_combout\,
	datac => \ConfigureCodec|ALT_INV_Selector11~0_combout\,
	datae => \ConfigureCodec|ALT_INV_R.BitCtr\(1),
	dataf => \ConfigureCodec|ALT_INV_Selector12~0_combout\,
	combout => \ConfigureCodec|Selector12~2_combout\);

-- Location: FF_X17_Y70_N19
\ConfigureCodec|R.BitCtr[1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \ConfigureCodec|Selector12~2_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ConfigureCodec|R.BitCtr\(1));

-- Location: LABCELL_X18_Y70_N24
\ConfigureCodec|NextR~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|NextR~9_combout\ = ( !\ConfigureCodec|R.BitCtr\(2) & ( (!\ConfigureCodec|R.BitCtr\(1) & !\ConfigureCodec|R.BitCtr[0]~DUPLICATE_q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1100000011000000110000001100000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ConfigureCodec|ALT_INV_R.BitCtr\(1),
	datac => \ConfigureCodec|ALT_INV_R.BitCtr[0]~DUPLICATE_q\,
	dataf => \ConfigureCodec|ALT_INV_R.BitCtr\(2),
	combout => \ConfigureCodec|NextR~9_combout\);

-- Location: LABCELL_X18_Y70_N30
\ConfigureCodec|Selector10~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Selector10~1_combout\ = ( \ConfigureCodec|Selector10~0_combout\ & ( \ConfigureCodec|NextStateAndOutput:vSclkFalling~0_combout\ & ( ((\ConfigureCodec|R.FrameState.Data1~q\ & (!\ConfigureCodec|R.BitCtr\(3) $ 
-- (!\ConfigureCodec|NextR~9_combout\)))) # (\ConfigureCodec|Selector5~0_combout\) ) ) ) # ( !\ConfigureCodec|Selector10~0_combout\ & ( \ConfigureCodec|NextStateAndOutput:vSclkFalling~0_combout\ & ( ((!\ConfigureCodec|R.BitCtr\(3) & 
-- (\ConfigureCodec|NextR~9_combout\ & \ConfigureCodec|R.FrameState.Data1~q\)) # (\ConfigureCodec|R.BitCtr\(3) & (!\ConfigureCodec|NextR~9_combout\))) # (\ConfigureCodec|Selector5~0_combout\) ) ) ) # ( !\ConfigureCodec|Selector10~0_combout\ & ( 
-- !\ConfigureCodec|NextStateAndOutput:vSclkFalling~0_combout\ & ( \ConfigureCodec|R.BitCtr\(3) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010101010101000000000000000001000110111111110000011011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ConfigureCodec|ALT_INV_R.BitCtr\(3),
	datab => \ConfigureCodec|ALT_INV_NextR~9_combout\,
	datac => \ConfigureCodec|ALT_INV_R.FrameState.Data1~q\,
	datad => \ConfigureCodec|ALT_INV_Selector5~0_combout\,
	datae => \ConfigureCodec|ALT_INV_Selector10~0_combout\,
	dataf => \ConfigureCodec|ALT_INV_NextStateAndOutput:vSclkFalling~0_combout\,
	combout => \ConfigureCodec|Selector10~1_combout\);

-- Location: LABCELL_X18_Y70_N48
\ConfigureCodec|Selector10~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Selector10~2_combout\ = ( \ConfigureCodec|R.BitCtr\(3) & ( \ConfigureCodec|R.FrameState.Data1~q\ & ( (((!\ConfigureCodec|Selector13~1_combout\) # (!\ConfigureCodec|NextStateAndOutput:vSclkFalling~0_combout\)) # 
-- (\ConfigureCodec|Selector10~1_combout\)) # (\ConfigureCodec|Selector1~0_combout\) ) ) ) # ( !\ConfigureCodec|R.BitCtr\(3) & ( \ConfigureCodec|R.FrameState.Data1~q\ & ( \ConfigureCodec|Selector10~1_combout\ ) ) ) # ( \ConfigureCodec|R.BitCtr\(3) & ( 
-- !\ConfigureCodec|R.FrameState.Data1~q\ & ( ((!\ConfigureCodec|Selector13~1_combout\) # (\ConfigureCodec|Selector10~1_combout\)) # (\ConfigureCodec|Selector1~0_combout\) ) ) ) # ( !\ConfigureCodec|R.BitCtr\(3) & ( !\ConfigureCodec|R.FrameState.Data1~q\ & ( 
-- \ConfigureCodec|Selector10~1_combout\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001100110011111101111111011100110011001100111111111111110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ConfigureCodec|ALT_INV_Selector1~0_combout\,
	datab => \ConfigureCodec|ALT_INV_Selector10~1_combout\,
	datac => \ConfigureCodec|ALT_INV_Selector13~1_combout\,
	datad => \ConfigureCodec|ALT_INV_NextStateAndOutput:vSclkFalling~0_combout\,
	datae => \ConfigureCodec|ALT_INV_R.BitCtr\(3),
	dataf => \ConfigureCodec|ALT_INV_R.FrameState.Data1~q\,
	combout => \ConfigureCodec|Selector10~2_combout\);

-- Location: FF_X18_Y70_N50
\ConfigureCodec|R.BitCtr[3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \ConfigureCodec|Selector10~2_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ConfigureCodec|R.BitCtr\(3));

-- Location: LABCELL_X18_Y70_N39
\ConfigureCodec|Selector6~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Selector6~0_combout\ = ( \ConfigureCodec|NextR~9_combout\ & ( (!\ConfigureCodec|NextStateAndOutput:vSclkFalling~0_combout\ & (((\ConfigureCodec|R.FrameState.Ack2~q\)))) # (\ConfigureCodec|NextStateAndOutput:vSclkFalling~0_combout\ & 
-- (\ConfigureCodec|R.BitCtr\(3) & (\ConfigureCodec|R.FrameState.Data1~q\))) ) ) # ( !\ConfigureCodec|NextR~9_combout\ & ( (!\ConfigureCodec|NextStateAndOutput:vSclkFalling~0_combout\ & \ConfigureCodec|R.FrameState.Ack2~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011001100000000001100110000000001110011010000000111001101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ConfigureCodec|ALT_INV_R.BitCtr\(3),
	datab => \ConfigureCodec|ALT_INV_NextStateAndOutput:vSclkFalling~0_combout\,
	datac => \ConfigureCodec|ALT_INV_R.FrameState.Data1~q\,
	datad => \ConfigureCodec|ALT_INV_R.FrameState.Ack2~q\,
	dataf => \ConfigureCodec|ALT_INV_NextR~9_combout\,
	combout => \ConfigureCodec|Selector6~0_combout\);

-- Location: FF_X18_Y70_N40
\ConfigureCodec|R.FrameState.Ack2\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \ConfigureCodec|Selector6~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ConfigureCodec|R.FrameState.Ack2~q\);

-- Location: LABCELL_X19_Y70_N54
\ConfigureCodec|Selector9~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Selector9~0_combout\ = ( \ConfigureCodec|R.FrameState.Stop~q\ & ( \ConfigureCodec|R.FrameState.Ack3~q\ ) ) # ( !\ConfigureCodec|R.FrameState.Stop~q\ & ( \ConfigureCodec|R.FrameState.Ack3~q\ & ( 
-- \ConfigureCodec|NextStateAndOutput:vSclkFalling~0_combout\ ) ) ) # ( \ConfigureCodec|R.FrameState.Stop~q\ & ( !\ConfigureCodec|R.FrameState.Ack3~q\ & ( (!\ConfigureCodec|NextStateAndOutput:vSclkFalling~0_combout\) # ((\ConfigureCodec|R.AckError~q\ & 
-- ((\ConfigureCodec|R.FrameState.Ack1~q\) # (\ConfigureCodec|R.FrameState.Ack2~q\)))) ) ) ) # ( !\ConfigureCodec|R.FrameState.Stop~q\ & ( !\ConfigureCodec|R.FrameState.Ack3~q\ & ( (\ConfigureCodec|R.AckError~q\ & 
-- (\ConfigureCodec|NextStateAndOutput:vSclkFalling~0_combout\ & ((\ConfigureCodec|R.FrameState.Ack1~q\) # (\ConfigureCodec|R.FrameState.Ack2~q\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000111111111110000011100000000111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ConfigureCodec|ALT_INV_R.FrameState.Ack2~q\,
	datab => \ConfigureCodec|ALT_INV_R.FrameState.Ack1~q\,
	datac => \ConfigureCodec|ALT_INV_R.AckError~q\,
	datad => \ConfigureCodec|ALT_INV_NextStateAndOutput:vSclkFalling~0_combout\,
	datae => \ConfigureCodec|ALT_INV_R.FrameState.Stop~q\,
	dataf => \ConfigureCodec|ALT_INV_R.FrameState.Ack3~q\,
	combout => \ConfigureCodec|Selector9~0_combout\);

-- Location: FF_X19_Y70_N56
\ConfigureCodec|R.FrameState.Stop\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \ConfigureCodec|Selector9~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ConfigureCodec|R.FrameState.Stop~q\);

-- Location: LABCELL_X19_Y70_N0
\ConfigureCodec|R.AddrCtr[6]~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|R.AddrCtr[6]~1_combout\ = ( !\ConfigureCodec|R.AckError~q\ & ( (\ConfigureCodec|R.FrameState.Stop~q\ & (!\ConfigureCodec|R.Sclk~q\ & \ConfigureCodec|R.Activity~q\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001010000000000000101000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ConfigureCodec|ALT_INV_R.FrameState.Stop~q\,
	datac => \ConfigureCodec|ALT_INV_R.Sclk~q\,
	datad => \ConfigureCodec|ALT_INV_R.Activity~q\,
	dataf => \ConfigureCodec|ALT_INV_R.AckError~q\,
	combout => \ConfigureCodec|R.AddrCtr[6]~1_combout\);

-- Location: LABCELL_X19_Y66_N6
\ConfigureCodec|R.Configured~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|R.Configured~0_combout\ = ( \ConfigureCodec|R.Configured~q\ & ( \GenStrobeI2C|oStrobe~q\ & ( (!\ConfigureCodec|R.AddrCtr[6]~0_combout\) # ((\ConfigureCodec|Equal0~1_combout\ & (\ConfigureCodec|Equal0~0_combout\ & 
-- \ConfigureCodec|R.AddrCtr[6]~1_combout\))) ) ) ) # ( !\ConfigureCodec|R.Configured~q\ & ( \GenStrobeI2C|oStrobe~q\ & ( (\ConfigureCodec|Equal0~1_combout\ & (\ConfigureCodec|Equal0~0_combout\ & \ConfigureCodec|R.AddrCtr[6]~1_combout\)) ) ) ) # ( 
-- \ConfigureCodec|R.Configured~q\ & ( !\GenStrobeI2C|oStrobe~q\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000111010101010101011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ConfigureCodec|ALT_INV_R.AddrCtr[6]~0_combout\,
	datab => \ConfigureCodec|ALT_INV_Equal0~1_combout\,
	datac => \ConfigureCodec|ALT_INV_Equal0~0_combout\,
	datad => \ConfigureCodec|ALT_INV_R.AddrCtr[6]~1_combout\,
	datae => \ConfigureCodec|ALT_INV_R.Configured~q\,
	dataf => \GenStrobeI2C|ALT_INV_oStrobe~q\,
	combout => \ConfigureCodec|R.Configured~0_combout\);

-- Location: FF_X19_Y66_N8
\ConfigureCodec|R.Configured\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \ConfigureCodec|R.Configured~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ConfigureCodec|R.Configured~q\);

-- Location: FF_X19_Y66_N35
\WaitCtr[0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \WaitCtr[0]~1_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => WaitCtr(0));

-- Location: LABCELL_X19_Y66_N48
\WaitCtr[1]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \WaitCtr[1]~0_combout\ = ( WaitCtr(1) & ( \GenStrobeI2C|oStrobe~q\ ) ) # ( !WaitCtr(1) & ( \GenStrobeI2C|oStrobe~q\ & ( (!\ConfigureCodec|R.Configured~q\ & WaitCtr(0)) ) ) ) # ( WaitCtr(1) & ( !\GenStrobeI2C|oStrobe~q\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100001100000011001111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ConfigureCodec|ALT_INV_R.Configured~q\,
	datac => ALT_INV_WaitCtr(0),
	datae => ALT_INV_WaitCtr(1),
	dataf => \GenStrobeI2C|ALT_INV_oStrobe~q\,
	combout => \WaitCtr[1]~0_combout\);

-- Location: FF_X19_Y66_N50
\WaitCtr[1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \WaitCtr[1]~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => WaitCtr(1));

-- Location: LABCELL_X19_Y66_N33
\WaitCtr[0]~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \WaitCtr[0]~1_combout\ = ( WaitCtr(0) & ( \GenStrobeI2C|oStrobe~q\ & ( (WaitCtr(1)) # (\ConfigureCodec|R.Configured~q\) ) ) ) # ( !WaitCtr(0) & ( \GenStrobeI2C|oStrobe~q\ & ( !\ConfigureCodec|R.Configured~q\ ) ) ) # ( WaitCtr(0) & ( 
-- !\GenStrobeI2C|oStrobe~q\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111111001100110011000011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ConfigureCodec|ALT_INV_R.Configured~q\,
	datad => ALT_INV_WaitCtr(1),
	datae => ALT_INV_WaitCtr(0),
	dataf => \GenStrobeI2C|ALT_INV_oStrobe~q\,
	combout => \WaitCtr[0]~1_combout\);

-- Location: FF_X19_Y66_N34
\WaitCtr[0]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \WaitCtr[0]~1_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \WaitCtr[0]~DUPLICATE_q\);

-- Location: LABCELL_X19_Y66_N27
\Start~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \Start~0_combout\ = ( \Start~q\ & ( \GenStrobeI2C|oStrobe~q\ & ( (\WaitCtr[0]~DUPLICATE_q\ & (!\ConfigureCodec|R.Configured~q\ & WaitCtr(1))) ) ) ) # ( !\Start~q\ & ( \GenStrobeI2C|oStrobe~q\ & ( (\WaitCtr[0]~DUPLICATE_q\ & 
-- (!\ConfigureCodec|R.Configured~q\ & WaitCtr(1))) ) ) ) # ( \Start~q\ & ( !\GenStrobeI2C|oStrobe~q\ & ( !\ConfigureCodec|R.Configured~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000010100000000000001010000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_WaitCtr[0]~DUPLICATE_q\,
	datac => \ConfigureCodec|ALT_INV_R.Configured~q\,
	datad => ALT_INV_WaitCtr(1),
	datae => \ALT_INV_Start~q\,
	dataf => \GenStrobeI2C|ALT_INV_oStrobe~q\,
	combout => \Start~0_combout\);

-- Location: FF_X19_Y66_N28
Start : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \Start~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \Start~q\);

-- Location: LABCELL_X19_Y66_N36
\ConfigureCodec|R.AddrCtr[6]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|R.AddrCtr[6]~0_combout\ = ( !\ConfigureCodec|R.Activity~q\ & ( \Start~q\ & ( !\ConfigureCodec|R.FrameState.Idle~DUPLICATE_q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011110000111100000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ConfigureCodec|ALT_INV_R.FrameState.Idle~DUPLICATE_q\,
	datae => \ConfigureCodec|ALT_INV_R.Activity~q\,
	dataf => \ALT_INV_Start~q\,
	combout => \ConfigureCodec|R.AddrCtr[6]~0_combout\);

-- Location: LABCELL_X19_Y66_N42
\ConfigureCodec|R.AddrCtr[6]~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|R.AddrCtr[6]~2_combout\ = ( \ConfigureCodec|Equal0~1_combout\ & ( (\GenStrobeI2C|oStrobe~q\ & (((!\ConfigureCodec|Equal0~0_combout\ & \ConfigureCodec|R.AddrCtr[6]~1_combout\)) # (\ConfigureCodec|R.AddrCtr[6]~0_combout\))) ) ) # ( 
-- !\ConfigureCodec|Equal0~1_combout\ & ( (\GenStrobeI2C|oStrobe~q\ & ((\ConfigureCodec|R.AddrCtr[6]~1_combout\) # (\ConfigureCodec|R.AddrCtr[6]~0_combout\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000100110011000100010011000100010001001100110001000100110001",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ConfigureCodec|ALT_INV_R.AddrCtr[6]~0_combout\,
	datab => \GenStrobeI2C|ALT_INV_oStrobe~q\,
	datac => \ConfigureCodec|ALT_INV_Equal0~0_combout\,
	datad => \ConfigureCodec|ALT_INV_R.AddrCtr[6]~1_combout\,
	datae => \ConfigureCodec|ALT_INV_Equal0~1_combout\,
	combout => \ConfigureCodec|R.AddrCtr[6]~2_combout\);

-- Location: FF_X21_Y70_N7
\ConfigureCodec|R.AddrCtr[2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \ConfigureCodec|Add0~1_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \ConfigureCodec|ALT_INV_R.Activity~q\,
	ena => \ConfigureCodec|R.AddrCtr[6]~2_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ConfigureCodec|R.AddrCtr\(2));

-- Location: FF_X21_Y70_N8
\ConfigureCodec|R.AddrCtr[2]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \ConfigureCodec|Add0~1_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \ConfigureCodec|ALT_INV_R.Activity~q\,
	ena => \ConfigureCodec|R.AddrCtr[6]~2_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ConfigureCodec|R.AddrCtr[2]~DUPLICATE_q\);

-- Location: FF_X21_Y70_N4
\ConfigureCodec|R.AddrCtr[1]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \ConfigureCodec|Add0~5_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \ConfigureCodec|ALT_INV_R.Activity~q\,
	ena => \ConfigureCodec|R.AddrCtr[6]~2_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ConfigureCodec|R.AddrCtr[1]~DUPLICATE_q\);

-- Location: LABCELL_X19_Y66_N0
\ConfigureCodec|Equal0~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Equal0~0_combout\ = ( !\ConfigureCodec|R.AddrCtr[2]~DUPLICATE_q\ & ( !\ConfigureCodec|R.AddrCtr[1]~DUPLICATE_q\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111111111111000000000000000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datae => \ConfigureCodec|ALT_INV_R.AddrCtr[2]~DUPLICATE_q\,
	dataf => \ConfigureCodec|ALT_INV_R.AddrCtr[1]~DUPLICATE_q\,
	combout => \ConfigureCodec|Equal0~0_combout\);

-- Location: LABCELL_X19_Y70_N3
\ConfigureCodec|R.Activity~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|R.Activity~0_combout\ = ( !\ConfigureCodec|R.Sclk~q\ & ( (\ConfigureCodec|R.FrameState.Stop~q\ & \GenStrobeI2C|oStrobe~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001010101000000000101010100000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ConfigureCodec|ALT_INV_R.FrameState.Stop~q\,
	datad => \GenStrobeI2C|ALT_INV_oStrobe~q\,
	dataf => \ConfigureCodec|ALT_INV_R.Sclk~q\,
	combout => \ConfigureCodec|R.Activity~0_combout\);

-- Location: LABCELL_X19_Y66_N15
\ConfigureCodec|Selector16~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Selector16~0_combout\ = ( !\ConfigureCodec|R.Activity~q\ & ( (!\ConfigureCodec|R.FrameState.Idle~DUPLICATE_q\ & (\Start~q\ & \GenStrobeI2C|oStrobe~q\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001000000010000000000000000000000010000000100000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ConfigureCodec|ALT_INV_R.FrameState.Idle~DUPLICATE_q\,
	datab => \ALT_INV_Start~q\,
	datac => \GenStrobeI2C|ALT_INV_oStrobe~q\,
	datae => \ConfigureCodec|ALT_INV_R.Activity~q\,
	combout => \ConfigureCodec|Selector16~0_combout\);

-- Location: LABCELL_X19_Y66_N54
\ConfigureCodec|R.Activity~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|R.Activity~1_combout\ = ( \ConfigureCodec|R.Activity~q\ & ( \ConfigureCodec|Selector16~0_combout\ ) ) # ( !\ConfigureCodec|R.Activity~q\ & ( \ConfigureCodec|Selector16~0_combout\ ) ) # ( \ConfigureCodec|R.Activity~q\ & ( 
-- !\ConfigureCodec|Selector16~0_combout\ & ( (!\ConfigureCodec|R.Activity~0_combout\) # ((!\ConfigureCodec|R.AckError~q\ & ((!\ConfigureCodec|Equal0~0_combout\) # (!\ConfigureCodec|Equal0~1_combout\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111101111000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ConfigureCodec|ALT_INV_Equal0~0_combout\,
	datab => \ConfigureCodec|ALT_INV_Equal0~1_combout\,
	datac => \ConfigureCodec|ALT_INV_R.Activity~0_combout\,
	datad => \ConfigureCodec|ALT_INV_R.AckError~q\,
	datae => \ConfigureCodec|ALT_INV_R.Activity~q\,
	dataf => \ConfigureCodec|ALT_INV_Selector16~0_combout\,
	combout => \ConfigureCodec|R.Activity~1_combout\);

-- Location: FF_X19_Y66_N56
\ConfigureCodec|R.Activity\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \ConfigureCodec|R.Activity~1_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ConfigureCodec|R.Activity~q\);

-- Location: LABCELL_X19_Y70_N12
\ConfigureCodec|Selector0~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Selector0~0_combout\ = ( \ConfigureCodec|R.Sclk~q\ & ( ((\GenStrobeI2C|oStrobe~q\ & \ConfigureCodec|R.Activity~q\)) # (\ConfigureCodec|R.FrameState.Idle~q\) ) ) # ( !\ConfigureCodec|R.Sclk~q\ & ( (!\GenStrobeI2C|oStrobe~q\ & 
-- (((\ConfigureCodec|R.FrameState.Idle~q\)))) # (\GenStrobeI2C|oStrobe~q\ & (!\ConfigureCodec|R.FrameState.Stop~q\ & ((\ConfigureCodec|R.FrameState.Idle~q\) # (\ConfigureCodec|R.Activity~q\)))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000011111010000100001111101000010001111111110001000111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \GenStrobeI2C|ALT_INV_oStrobe~q\,
	datab => \ConfigureCodec|ALT_INV_R.Activity~q\,
	datac => \ConfigureCodec|ALT_INV_R.FrameState.Stop~q\,
	datad => \ConfigureCodec|ALT_INV_R.FrameState.Idle~q\,
	dataf => \ConfigureCodec|ALT_INV_R.Sclk~q\,
	combout => \ConfigureCodec|Selector0~0_combout\);

-- Location: FF_X19_Y70_N14
\ConfigureCodec|R.FrameState.Idle\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \ConfigureCodec|Selector0~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ConfigureCodec|R.FrameState.Idle~q\);

-- Location: LABCELL_X19_Y70_N18
\ConfigureCodec|Selector14~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Selector14~0_combout\ = ( \ConfigureCodec|R.Activity~q\ & ( (!\GenStrobeI2C|oStrobe~q\ & (((\ConfigureCodec|R.Sclk~q\)))) # (\GenStrobeI2C|oStrobe~q\ & (\ConfigureCodec|R.FrameState.Idle~q\ & (!\ConfigureCodec|R.FrameState.Stop~q\ & 
-- !\ConfigureCodec|R.Sclk~q\))) ) ) # ( !\ConfigureCodec|R.Activity~q\ & ( \ConfigureCodec|R.Sclk~q\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011111111000000001111111100010000101010100001000010101010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \GenStrobeI2C|ALT_INV_oStrobe~q\,
	datab => \ConfigureCodec|ALT_INV_R.FrameState.Idle~q\,
	datac => \ConfigureCodec|ALT_INV_R.FrameState.Stop~q\,
	datad => \ConfigureCodec|ALT_INV_R.Sclk~q\,
	dataf => \ConfigureCodec|ALT_INV_R.Activity~q\,
	combout => \ConfigureCodec|Selector14~0_combout\);

-- Location: FF_X19_Y70_N19
\ConfigureCodec|R.Sclk\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \ConfigureCodec|Selector14~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ConfigureCodec|R.Sclk~q\);

-- Location: LABCELL_X19_Y70_N15
\ConfigureCodec|Selector15~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Selector15~1_combout\ = ( \ConfigureCodec|R.FrameState.Idle~q\ & ( !\ConfigureCodec|R.FrameState.Start~q\ ) ) # ( !\ConfigureCodec|R.FrameState.Idle~q\ & ( (\ConfigureCodec|R.Activity~q\ & (!\ConfigureCodec|R.FrameState.Start~q\ & 
-- \GenStrobeI2C|oStrobe~q\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000110000000000000011000011110000111100001111000011110000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ConfigureCodec|ALT_INV_R.Activity~q\,
	datac => \ConfigureCodec|ALT_INV_R.FrameState.Start~q\,
	datad => \GenStrobeI2C|ALT_INV_oStrobe~q\,
	dataf => \ConfigureCodec|ALT_INV_R.FrameState.Idle~q\,
	combout => \ConfigureCodec|Selector15~1_combout\);

-- Location: LABCELL_X18_Y70_N12
\ConfigureCodec|Selector15~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Selector15~2_combout\ = ( \ConfigureCodec|Selector13~0_combout\ & ( (!\ConfigureCodec|R.Activity~0_combout\ & ((\ConfigureCodec|R.Sdin~q\) # (\ConfigureCodec|Selector15~1_combout\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000001010000111100000101000011110000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ConfigureCodec|ALT_INV_Selector15~1_combout\,
	datac => \ConfigureCodec|ALT_INV_R.Activity~0_combout\,
	datad => \ConfigureCodec|ALT_INV_R.Sdin~q\,
	dataf => \ConfigureCodec|ALT_INV_Selector13~0_combout\,
	combout => \ConfigureCodec|Selector15~2_combout\);

-- Location: LABCELL_X19_Y70_N24
\ConfigureCodec|R.Data[15]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|R.Data[15]~0_combout\ = (\GenStrobeI2C|oStrobe~q\ & (\ConfigureCodec|R.FrameState.Start~q\ & \ConfigureCodec|R.Activity~q\))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000010001000000000001000100000000000100010000000000010001",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \GenStrobeI2C|ALT_INV_oStrobe~q\,
	datab => \ConfigureCodec|ALT_INV_R.FrameState.Start~q\,
	datad => \ConfigureCodec|ALT_INV_R.Activity~q\,
	combout => \ConfigureCodec|R.Data[15]~0_combout\);

-- Location: FF_X18_Y70_N5
\ConfigureCodec|R.Data[11]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	asdata => \ConfigureCodec|R.AddrCtr[2]~DUPLICATE_q\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \ConfigureCodec|R.Data[15]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ConfigureCodec|R.Data\(11));

-- Location: MLABCELL_X21_Y70_N24
\ConfigureCodec|Mux0~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Mux0~0_combout\ = ( \ConfigureCodec|R.AddrCtr\(2) & ( (!\ConfigureCodec|R.AddrCtr\(1) & !\ConfigureCodec|R.AddrCtr\(0)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000010100000101000001010000010100000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ConfigureCodec|ALT_INV_R.AddrCtr\(1),
	datac => \ConfigureCodec|ALT_INV_R.AddrCtr\(0),
	dataf => \ConfigureCodec|ALT_INV_R.AddrCtr\(2),
	combout => \ConfigureCodec|Mux0~0_combout\);

-- Location: FF_X21_Y70_N25
\ConfigureCodec|R.Data[7]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \ConfigureCodec|Mux0~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	ena => \ConfigureCodec|R.Data[15]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ConfigureCodec|R.Data\(7));

-- Location: LABCELL_X18_Y70_N6
\ConfigureCodec|Mux4~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Mux4~0_combout\ = ( !\ConfigureCodec|R.AddrCtr\(3) & ( !\ConfigureCodec|R.AddrCtr[2]~DUPLICATE_q\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111000011110000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \ConfigureCodec|ALT_INV_R.AddrCtr[2]~DUPLICATE_q\,
	dataf => \ConfigureCodec|ALT_INV_R.AddrCtr\(3),
	combout => \ConfigureCodec|Mux4~0_combout\);

-- Location: FF_X18_Y70_N8
\ConfigureCodec|R.Data[3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \ConfigureCodec|Mux4~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	ena => \ConfigureCodec|R.Data[15]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ConfigureCodec|R.Data\(3));

-- Location: FF_X18_Y70_N20
\ConfigureCodec|R.Data[15]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	asdata => \ConfigureCodec|R.AddrCtr\(6),
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \ConfigureCodec|R.Data[15]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ConfigureCodec|R.Data\(15));

-- Location: LABCELL_X18_Y70_N18
\ConfigureCodec|Mux9~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Mux9~3_combout\ = ( \ConfigureCodec|R.Data\(15) & ( \ConfigureCodec|R.BitCtr\(3) & ( (\ConfigureCodec|R.BitCtr\(2)) # (\ConfigureCodec|R.Data\(11)) ) ) ) # ( !\ConfigureCodec|R.Data\(15) & ( \ConfigureCodec|R.BitCtr\(3) & ( 
-- (\ConfigureCodec|R.Data\(11) & !\ConfigureCodec|R.BitCtr\(2)) ) ) ) # ( \ConfigureCodec|R.Data\(15) & ( !\ConfigureCodec|R.BitCtr\(3) & ( (!\ConfigureCodec|R.BitCtr\(2) & ((\ConfigureCodec|R.Data\(3)))) # (\ConfigureCodec|R.BitCtr\(2) & 
-- (\ConfigureCodec|R.Data\(7))) ) ) ) # ( !\ConfigureCodec|R.Data\(15) & ( !\ConfigureCodec|R.BitCtr\(3) & ( (!\ConfigureCodec|R.BitCtr\(2) & ((\ConfigureCodec|R.Data\(3)))) # (\ConfigureCodec|R.BitCtr\(2) & (\ConfigureCodec|R.Data\(7))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001111001111000000111100111101000100010001000111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ConfigureCodec|ALT_INV_R.Data\(11),
	datab => \ConfigureCodec|ALT_INV_R.BitCtr\(2),
	datac => \ConfigureCodec|ALT_INV_R.Data\(7),
	datad => \ConfigureCodec|ALT_INV_R.Data\(3),
	datae => \ConfigureCodec|ALT_INV_R.Data\(15),
	dataf => \ConfigureCodec|ALT_INV_R.BitCtr\(3),
	combout => \ConfigureCodec|Mux9~3_combout\);

-- Location: MLABCELL_X21_Y70_N36
\ConfigureCodec|Mux6~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Mux6~0_combout\ = ( \ConfigureCodec|R.AddrCtr\(2) & ( (!\ConfigureCodec|R.AddrCtr\(3) & ((!\ConfigureCodec|R.AddrCtr\(0)) # (\ConfigureCodec|R.AddrCtr\(1)))) ) ) # ( !\ConfigureCodec|R.AddrCtr\(2) & ( (!\ConfigureCodec|R.AddrCtr\(1) & 
-- ((!\ConfigureCodec|R.AddrCtr\(0)) # (!\ConfigureCodec|R.AddrCtr\(3)))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1110000011100000111000001110000010001100100011001000110010001100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ConfigureCodec|ALT_INV_R.AddrCtr\(0),
	datab => \ConfigureCodec|ALT_INV_R.AddrCtr\(3),
	datac => \ConfigureCodec|ALT_INV_R.AddrCtr\(1),
	dataf => \ConfigureCodec|ALT_INV_R.AddrCtr\(2),
	combout => \ConfigureCodec|Mux6~0_combout\);

-- Location: FF_X21_Y70_N38
\ConfigureCodec|R.Data[1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \ConfigureCodec|Mux6~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	ena => \ConfigureCodec|R.Data[15]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ConfigureCodec|R.Data\(1));

-- Location: FF_X21_Y70_N59
\ConfigureCodec|R.Data[9]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	asdata => \ConfigureCodec|R.AddrCtr\(0),
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \ConfigureCodec|R.Data[15]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ConfigureCodec|R.Data\(9));

-- Location: FF_X21_Y70_N56
\ConfigureCodec|R.Data[13]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	asdata => \ConfigureCodec|R.AddrCtr\(4),
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \ConfigureCodec|R.Data[15]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ConfigureCodec|R.Data\(13));

-- Location: MLABCELL_X21_Y70_N39
\ConfigureCodec|Mux2~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Mux2~0_combout\ = ( \ConfigureCodec|R.AddrCtr\(2) & ( (!\ConfigureCodec|R.AddrCtr\(0) & (!\ConfigureCodec|R.AddrCtr\(3) & \ConfigureCodec|R.AddrCtr\(1))) ) ) # ( !\ConfigureCodec|R.AddrCtr\(2) & ( (!\ConfigureCodec|R.AddrCtr\(3) & 
-- ((\ConfigureCodec|R.AddrCtr\(1)))) # (\ConfigureCodec|R.AddrCtr\(3) & (!\ConfigureCodec|R.AddrCtr\(0) & !\ConfigureCodec|R.AddrCtr\(1))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000101011110000000010101111000000000000101000000000000010100000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ConfigureCodec|ALT_INV_R.AddrCtr\(0),
	datac => \ConfigureCodec|ALT_INV_R.AddrCtr\(3),
	datad => \ConfigureCodec|ALT_INV_R.AddrCtr\(1),
	dataf => \ConfigureCodec|ALT_INV_R.AddrCtr\(2),
	combout => \ConfigureCodec|Mux2~0_combout\);

-- Location: FF_X21_Y70_N41
\ConfigureCodec|R.Data[5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \ConfigureCodec|Mux2~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	ena => \ConfigureCodec|R.Data[15]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ConfigureCodec|R.Data\(5));

-- Location: MLABCELL_X21_Y70_N54
\ConfigureCodec|Mux9~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Mux9~2_combout\ = ( \ConfigureCodec|R.Data\(13) & ( \ConfigureCodec|R.Data\(5) & ( ((!\ConfigureCodec|R.BitCtr[3]~DUPLICATE_q\ & (\ConfigureCodec|R.Data\(1))) # (\ConfigureCodec|R.BitCtr[3]~DUPLICATE_q\ & ((\ConfigureCodec|R.Data\(9))))) # 
-- (\ConfigureCodec|R.BitCtr\(2)) ) ) ) # ( !\ConfigureCodec|R.Data\(13) & ( \ConfigureCodec|R.Data\(5) & ( (!\ConfigureCodec|R.BitCtr\(2) & ((!\ConfigureCodec|R.BitCtr[3]~DUPLICATE_q\ & (\ConfigureCodec|R.Data\(1))) # 
-- (\ConfigureCodec|R.BitCtr[3]~DUPLICATE_q\ & ((\ConfigureCodec|R.Data\(9)))))) # (\ConfigureCodec|R.BitCtr\(2) & (!\ConfigureCodec|R.BitCtr[3]~DUPLICATE_q\)) ) ) ) # ( \ConfigureCodec|R.Data\(13) & ( !\ConfigureCodec|R.Data\(5) & ( 
-- (!\ConfigureCodec|R.BitCtr\(2) & ((!\ConfigureCodec|R.BitCtr[3]~DUPLICATE_q\ & (\ConfigureCodec|R.Data\(1))) # (\ConfigureCodec|R.BitCtr[3]~DUPLICATE_q\ & ((\ConfigureCodec|R.Data\(9)))))) # (\ConfigureCodec|R.BitCtr\(2) & 
-- (\ConfigureCodec|R.BitCtr[3]~DUPLICATE_q\)) ) ) ) # ( !\ConfigureCodec|R.Data\(13) & ( !\ConfigureCodec|R.Data\(5) & ( (!\ConfigureCodec|R.BitCtr\(2) & ((!\ConfigureCodec|R.BitCtr[3]~DUPLICATE_q\ & (\ConfigureCodec|R.Data\(1))) # 
-- (\ConfigureCodec|R.BitCtr[3]~DUPLICATE_q\ & ((\ConfigureCodec|R.Data\(9)))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000100000101010000110010011101101001100011011100101110101111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ConfigureCodec|ALT_INV_R.BitCtr\(2),
	datab => \ConfigureCodec|ALT_INV_R.BitCtr[3]~DUPLICATE_q\,
	datac => \ConfigureCodec|ALT_INV_R.Data\(1),
	datad => \ConfigureCodec|ALT_INV_R.Data\(9),
	datae => \ConfigureCodec|ALT_INV_R.Data\(13),
	dataf => \ConfigureCodec|ALT_INV_R.Data\(5),
	combout => \ConfigureCodec|Mux9~2_combout\);

-- Location: MLABCELL_X21_Y70_N27
\ConfigureCodec|Mux5~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Mux5~0_combout\ = ( !\ConfigureCodec|R.AddrCtr\(2) & ( (!\ConfigureCodec|R.AddrCtr\(1) & !\ConfigureCodec|R.AddrCtr\(3)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1010000010100000101000001010000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ConfigureCodec|ALT_INV_R.AddrCtr\(1),
	datac => \ConfigureCodec|ALT_INV_R.AddrCtr\(3),
	dataf => \ConfigureCodec|ALT_INV_R.AddrCtr\(2),
	combout => \ConfigureCodec|Mux5~0_combout\);

-- Location: FF_X21_Y70_N29
\ConfigureCodec|R.Data[2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \ConfigureCodec|Mux5~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	ena => \ConfigureCodec|R.Data[15]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ConfigureCodec|R.Data\(2));

-- Location: FF_X21_Y70_N47
\ConfigureCodec|R.Data[14]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	asdata => \ConfigureCodec|R.AddrCtr\(5),
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \ConfigureCodec|R.Data[15]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ConfigureCodec|R.Data\(14));

-- Location: FF_X21_Y70_N44
\ConfigureCodec|R.Data[10]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	asdata => \ConfigureCodec|R.AddrCtr\(1),
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \ConfigureCodec|R.Data[15]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ConfigureCodec|R.Data\(10));

-- Location: MLABCELL_X21_Y70_N33
\ConfigureCodec|Mux1~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Mux1~0_combout\ = ( \ConfigureCodec|R.AddrCtr\(2) & ( !\ConfigureCodec|R.AddrCtr\(0) ) ) # ( !\ConfigureCodec|R.AddrCtr\(2) & ( \ConfigureCodec|R.AddrCtr\(1) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011111111000000001111111110101010101010101010101010101010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ConfigureCodec|ALT_INV_R.AddrCtr\(0),
	datad => \ConfigureCodec|ALT_INV_R.AddrCtr\(1),
	dataf => \ConfigureCodec|ALT_INV_R.AddrCtr\(2),
	combout => \ConfigureCodec|Mux1~0_combout\);

-- Location: FF_X21_Y70_N35
\ConfigureCodec|R.Data[6]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \ConfigureCodec|Mux1~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	ena => \ConfigureCodec|R.Data[15]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ConfigureCodec|R.Data\(6));

-- Location: MLABCELL_X21_Y70_N42
\ConfigureCodec|Mux9~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Mux9~1_combout\ = ( \ConfigureCodec|R.Data\(10) & ( \ConfigureCodec|R.Data\(6) & ( (!\ConfigureCodec|R.BitCtr\(2) & (((\ConfigureCodec|R.BitCtr[3]~DUPLICATE_q\)) # (\ConfigureCodec|R.Data\(2)))) # (\ConfigureCodec|R.BitCtr\(2) & 
-- (((!\ConfigureCodec|R.BitCtr[3]~DUPLICATE_q\) # (\ConfigureCodec|R.Data\(14))))) ) ) ) # ( !\ConfigureCodec|R.Data\(10) & ( \ConfigureCodec|R.Data\(6) & ( (!\ConfigureCodec|R.BitCtr\(2) & (\ConfigureCodec|R.Data\(2) & 
-- ((!\ConfigureCodec|R.BitCtr[3]~DUPLICATE_q\)))) # (\ConfigureCodec|R.BitCtr\(2) & (((!\ConfigureCodec|R.BitCtr[3]~DUPLICATE_q\) # (\ConfigureCodec|R.Data\(14))))) ) ) ) # ( \ConfigureCodec|R.Data\(10) & ( !\ConfigureCodec|R.Data\(6) & ( 
-- (!\ConfigureCodec|R.BitCtr\(2) & (((\ConfigureCodec|R.BitCtr[3]~DUPLICATE_q\)) # (\ConfigureCodec|R.Data\(2)))) # (\ConfigureCodec|R.BitCtr\(2) & (((\ConfigureCodec|R.Data\(14) & \ConfigureCodec|R.BitCtr[3]~DUPLICATE_q\)))) ) ) ) # ( 
-- !\ConfigureCodec|R.Data\(10) & ( !\ConfigureCodec|R.Data\(6) & ( (!\ConfigureCodec|R.BitCtr\(2) & (\ConfigureCodec|R.Data\(2) & ((!\ConfigureCodec|R.BitCtr[3]~DUPLICATE_q\)))) # (\ConfigureCodec|R.BitCtr\(2) & (((\ConfigureCodec|R.Data\(14) & 
-- \ConfigureCodec|R.BitCtr[3]~DUPLICATE_q\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101000000000011010100001111001101011111000000110101111111110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ConfigureCodec|ALT_INV_R.Data\(2),
	datab => \ConfigureCodec|ALT_INV_R.Data\(14),
	datac => \ConfigureCodec|ALT_INV_R.BitCtr\(2),
	datad => \ConfigureCodec|ALT_INV_R.BitCtr[3]~DUPLICATE_q\,
	datae => \ConfigureCodec|ALT_INV_R.Data\(10),
	dataf => \ConfigureCodec|ALT_INV_R.Data\(6),
	combout => \ConfigureCodec|Mux9~1_combout\);

-- Location: MLABCELL_X21_Y70_N51
\ConfigureCodec|Mux3~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Mux3~0_combout\ = ( \ConfigureCodec|R.AddrCtr\(2) & ( (!\ConfigureCodec|R.AddrCtr\(0) & (!\ConfigureCodec|R.AddrCtr\(3) & !\ConfigureCodec|R.AddrCtr\(1))) ) ) # ( !\ConfigureCodec|R.AddrCtr\(2) & ( !\ConfigureCodec|R.AddrCtr\(3) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1100110011001100110011001100110010001000000000001000100000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ConfigureCodec|ALT_INV_R.AddrCtr\(0),
	datab => \ConfigureCodec|ALT_INV_R.AddrCtr\(3),
	datad => \ConfigureCodec|ALT_INV_R.AddrCtr\(1),
	dataf => \ConfigureCodec|ALT_INV_R.AddrCtr\(2),
	combout => \ConfigureCodec|Mux3~0_combout\);

-- Location: FF_X21_Y70_N52
\ConfigureCodec|R.Data[4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \ConfigureCodec|Mux3~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	ena => \ConfigureCodec|R.Data[15]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ConfigureCodec|R.Data\(4));

-- Location: FF_X18_Y70_N11
\ConfigureCodec|R.Data[12]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	asdata => \ConfigureCodec|R.AddrCtr\(3),
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \ConfigureCodec|R.Data[15]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ConfigureCodec|R.Data\(12));

-- Location: MLABCELL_X21_Y70_N30
\ConfigureCodec|Mux7~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Mux7~0_combout\ = ( \ConfigureCodec|R.AddrCtr\(2) & ( (\ConfigureCodec|R.AddrCtr\(0) & !\ConfigureCodec|R.AddrCtr\(1)) ) ) # ( !\ConfigureCodec|R.AddrCtr\(2) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111111111111111111111111111101010000010100000101000001010000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ConfigureCodec|ALT_INV_R.AddrCtr\(0),
	datac => \ConfigureCodec|ALT_INV_R.AddrCtr\(1),
	dataf => \ConfigureCodec|ALT_INV_R.AddrCtr\(2),
	combout => \ConfigureCodec|Mux7~0_combout\);

-- Location: FF_X21_Y70_N31
\ConfigureCodec|R.Data[0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \ConfigureCodec|Mux7~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	ena => \ConfigureCodec|R.Data[15]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ConfigureCodec|R.Data\(0));

-- Location: LABCELL_X18_Y70_N9
\ConfigureCodec|Mux9~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Mux9~0_combout\ = ( \ConfigureCodec|R.Data\(0) & ( (!\ConfigureCodec|R.BitCtr\(3) & ((!\ConfigureCodec|R.BitCtr\(2)) # ((\ConfigureCodec|R.Data\(4))))) # (\ConfigureCodec|R.BitCtr\(3) & (\ConfigureCodec|R.BitCtr\(2) & 
-- ((\ConfigureCodec|R.Data\(12))))) ) ) # ( !\ConfigureCodec|R.Data\(0) & ( (\ConfigureCodec|R.BitCtr\(2) & ((!\ConfigureCodec|R.BitCtr\(3) & (\ConfigureCodec|R.Data\(4))) # (\ConfigureCodec|R.BitCtr\(3) & ((\ConfigureCodec|R.Data\(12)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001000010011000000100001001110001010100110111000101010011011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ConfigureCodec|ALT_INV_R.BitCtr\(3),
	datab => \ConfigureCodec|ALT_INV_R.BitCtr\(2),
	datac => \ConfigureCodec|ALT_INV_R.Data\(4),
	datad => \ConfigureCodec|ALT_INV_R.Data\(12),
	dataf => \ConfigureCodec|ALT_INV_R.Data\(0),
	combout => \ConfigureCodec|Mux9~0_combout\);

-- Location: LABCELL_X18_Y70_N0
\ConfigureCodec|Mux9~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Mux9~4_combout\ = ( \ConfigureCodec|Mux9~1_combout\ & ( \ConfigureCodec|Mux9~0_combout\ & ( (!\ConfigureCodec|R.BitCtr[0]~DUPLICATE_q\) # ((!\ConfigureCodec|R.BitCtr\(1) & ((\ConfigureCodec|Mux9~2_combout\))) # 
-- (\ConfigureCodec|R.BitCtr\(1) & (\ConfigureCodec|Mux9~3_combout\))) ) ) ) # ( !\ConfigureCodec|Mux9~1_combout\ & ( \ConfigureCodec|Mux9~0_combout\ & ( (!\ConfigureCodec|R.BitCtr\(1) & (((!\ConfigureCodec|R.BitCtr[0]~DUPLICATE_q\) # 
-- (\ConfigureCodec|Mux9~2_combout\)))) # (\ConfigureCodec|R.BitCtr\(1) & (\ConfigureCodec|Mux9~3_combout\ & ((\ConfigureCodec|R.BitCtr[0]~DUPLICATE_q\)))) ) ) ) # ( \ConfigureCodec|Mux9~1_combout\ & ( !\ConfigureCodec|Mux9~0_combout\ & ( 
-- (!\ConfigureCodec|R.BitCtr\(1) & (((\ConfigureCodec|Mux9~2_combout\ & \ConfigureCodec|R.BitCtr[0]~DUPLICATE_q\)))) # (\ConfigureCodec|R.BitCtr\(1) & (((!\ConfigureCodec|R.BitCtr[0]~DUPLICATE_q\)) # (\ConfigureCodec|Mux9~3_combout\))) ) ) ) # ( 
-- !\ConfigureCodec|Mux9~1_combout\ & ( !\ConfigureCodec|Mux9~0_combout\ & ( (\ConfigureCodec|R.BitCtr[0]~DUPLICATE_q\ & ((!\ConfigureCodec|R.BitCtr\(1) & ((\ConfigureCodec|Mux9~2_combout\))) # (\ConfigureCodec|R.BitCtr\(1) & 
-- (\ConfigureCodec|Mux9~3_combout\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000011101001100110001110111001100000111011111111100011101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ConfigureCodec|ALT_INV_Mux9~3_combout\,
	datab => \ConfigureCodec|ALT_INV_R.BitCtr\(1),
	datac => \ConfigureCodec|ALT_INV_Mux9~2_combout\,
	datad => \ConfigureCodec|ALT_INV_R.BitCtr[0]~DUPLICATE_q\,
	datae => \ConfigureCodec|ALT_INV_Mux9~1_combout\,
	dataf => \ConfigureCodec|ALT_INV_Mux9~0_combout\,
	combout => \ConfigureCodec|Mux9~4_combout\);

-- Location: LABCELL_X18_Y70_N15
\ConfigureCodec|Selector15~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Selector15~0_combout\ = ( \ConfigureCodec|R.BitCtr\(2) & ( (!\ConfigureCodec|R.BitCtr[0]~DUPLICATE_q\ & (!\ConfigureCodec|R.BitCtr\(1) & \ConfigureCodec|R.FrameState.Address~q\)) ) ) # ( !\ConfigureCodec|R.BitCtr\(2) & ( 
-- (\ConfigureCodec|R.BitCtr[0]~DUPLICATE_q\ & \ConfigureCodec|R.FrameState.Address~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000110011000000000011001100000000110000000000000011000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \ConfigureCodec|ALT_INV_R.BitCtr[0]~DUPLICATE_q\,
	datac => \ConfigureCodec|ALT_INV_R.BitCtr\(1),
	datad => \ConfigureCodec|ALT_INV_R.FrameState.Address~q\,
	dataf => \ConfigureCodec|ALT_INV_R.BitCtr\(2),
	combout => \ConfigureCodec|Selector15~0_combout\);

-- Location: LABCELL_X18_Y70_N42
\ConfigureCodec|Selector15~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \ConfigureCodec|Selector15~3_combout\ = ( !\ConfigureCodec|Selector15~0_combout\ & ( (\ConfigureCodec|Selector15~2_combout\ & ((!\ConfigureCodec|Mux9~4_combout\) # ((!\ConfigureCodec|R.FrameState.Data1~q\ & !\ConfigureCodec|R.FrameState.Data2~q\)))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001100100000001100110010000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ConfigureCodec|ALT_INV_R.FrameState.Data1~q\,
	datab => \ConfigureCodec|ALT_INV_Selector15~2_combout\,
	datac => \ConfigureCodec|ALT_INV_R.FrameState.Data2~q\,
	datad => \ConfigureCodec|ALT_INV_Mux9~4_combout\,
	dataf => \ConfigureCodec|ALT_INV_Selector15~0_combout\,
	combout => \ConfigureCodec|Selector15~3_combout\);

-- Location: FF_X18_Y70_N43
\ConfigureCodec|R.Sdin\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \ConfigureCodec|Selector15~3_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ConfigureCodec|R.Sdin~q\);

-- Location: CLKCTRL_G4
\iClk~inputCLKENA0\ : cyclonev_clkena
-- pragma translate_off
GENERIC MAP (
	clock_type => "global clock",
	disable_mode => "low",
	ena_register_mode => "always enabled",
	ena_register_power_up => "high",
	test_syn => "high")
-- pragma translate_on
PORT MAP (
	inclk => \iClk~input_o\,
	outclk => \iClk~inputCLKENA0_outclk\);

-- Location: IOIBUF_X12_Y0_N18
\iSwitch[0]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_iSwitch(0),
	o => \iSwitch[0]~input_o\);

-- Location: DDIOINCELL_X12_Y0_N31
\SyncSwitchInput|Metastable[0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \iSwitch[0]~input_o\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \SyncSwitchInput|Metastable\(0));

-- Location: FF_X24_Y60_N50
\SyncSwitchInput|Metastable[1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	asdata => \SyncSwitchInput|Metastable\(0),
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \SyncSwitchInput|Metastable\(1));

-- Location: FF_X19_Y66_N7
\ConfigureCodec|R.Configured~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \ConfigureCodec|R.Configured~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \ConfigureCodec|R.Configured~DUPLICATE_q\);

-- Location: MLABCELL_X15_Y64_N30
\GenClks|Add0~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \GenClks|Add0~9_sumout\ = SUM(( \GenClks|BitCounter\(0) ) + ( VCC ) + ( !VCC ))
-- \GenClks|Add0~10\ = CARRY(( \GenClks|BitCounter\(0) ) + ( VCC ) + ( !VCC ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \GenClks|ALT_INV_BitCounter\(0),
	cin => GND,
	sumout => \GenClks|Add0~9_sumout\,
	cout => \GenClks|Add0~10\);

-- Location: MLABCELL_X15_Y64_N15
\GenClks|ClkCounter[0]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \GenClks|ClkCounter[0]~0_combout\ = ( !\GenClks|ClkCounter\(0) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111111111111000000000000000011111111111111110000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datae => \GenClks|ALT_INV_ClkCounter\(0),
	combout => \GenClks|ClkCounter[0]~0_combout\);

-- Location: FF_X15_Y64_N16
\GenClks|ClkCounter[0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \GenClks|ClkCounter[0]~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \GenClks|ClkCounter\(0));

-- Location: MLABCELL_X15_Y64_N0
\GenClks|BMclk~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \GenClks|BMclk~0_combout\ = ( !\GenClks|BMclk~q\ & ( \GenClks|ClkCounter\(0) ) ) # ( \GenClks|BMclk~q\ & ( !\GenClks|ClkCounter\(0) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111111111111111111110000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datae => \GenClks|ALT_INV_BMclk~q\,
	dataf => \GenClks|ALT_INV_ClkCounter\(0),
	combout => \GenClks|BMclk~0_combout\);

-- Location: FF_X15_Y64_N1
\GenClks|BMclk\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \GenClks|BMclk~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \GenClks|BMclk~q\);

-- Location: LABCELL_X13_Y64_N0
\GenClks|ADClrc~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \GenClks|ADClrc~0_combout\ = ( \GenClks|ClkCounter\(0) & ( \GenClks|BMclk~q\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000000000001111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datae => \GenClks|ALT_INV_ClkCounter\(0),
	dataf => \GenClks|ALT_INV_BMclk~q\,
	combout => \GenClks|ADClrc~0_combout\);

-- Location: FF_X15_Y64_N32
\GenClks|BitCounter[0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \GenClks|Add0~9_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	ena => \GenClks|ADClrc~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \GenClks|BitCounter\(0));

-- Location: MLABCELL_X15_Y64_N33
\GenClks|Add0~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \GenClks|Add0~5_sumout\ = SUM(( \GenClks|BitCounter\(1) ) + ( GND ) + ( \GenClks|Add0~10\ ))
-- \GenClks|Add0~6\ = CARRY(( \GenClks|BitCounter\(1) ) + ( GND ) + ( \GenClks|Add0~10\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \GenClks|ALT_INV_BitCounter\(1),
	cin => \GenClks|Add0~10\,
	sumout => \GenClks|Add0~5_sumout\,
	cout => \GenClks|Add0~6\);

-- Location: FF_X15_Y64_N35
\GenClks|BitCounter[1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \GenClks|Add0~5_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	ena => \GenClks|ADClrc~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \GenClks|BitCounter\(1));

-- Location: MLABCELL_X15_Y64_N36
\GenClks|Add0~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \GenClks|Add0~1_sumout\ = SUM(( \GenClks|BitCounter\(2) ) + ( GND ) + ( \GenClks|Add0~6\ ))
-- \GenClks|Add0~2\ = CARRY(( \GenClks|BitCounter\(2) ) + ( GND ) + ( \GenClks|Add0~6\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \GenClks|ALT_INV_BitCounter\(2),
	cin => \GenClks|Add0~6\,
	sumout => \GenClks|Add0~1_sumout\,
	cout => \GenClks|Add0~2\);

-- Location: FF_X15_Y64_N38
\GenClks|BitCounter[2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \GenClks|Add0~1_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	ena => \GenClks|ADClrc~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \GenClks|BitCounter\(2));

-- Location: MLABCELL_X15_Y64_N39
\GenClks|Add0~29\ : cyclonev_lcell_comb
-- Equation(s):
-- \GenClks|Add0~29_sumout\ = SUM(( \GenClks|BitCounter\(3) ) + ( GND ) + ( \GenClks|Add0~2\ ))
-- \GenClks|Add0~30\ = CARRY(( \GenClks|BitCounter\(3) ) + ( GND ) + ( \GenClks|Add0~2\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \GenClks|ALT_INV_BitCounter\(3),
	cin => \GenClks|Add0~2\,
	sumout => \GenClks|Add0~29_sumout\,
	cout => \GenClks|Add0~30\);

-- Location: FF_X15_Y64_N34
\GenClks|BitCounter[1]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \GenClks|Add0~5_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	ena => \GenClks|ADClrc~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \GenClks|BitCounter[1]~DUPLICATE_q\);

-- Location: MLABCELL_X15_Y64_N9
\GenClks|BitCounter~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \GenClks|BitCounter~1_combout\ = ( \GenClks|Equal0~0_combout\ & ( (\GenClks|Add0~29_sumout\ & ((!\GenClks|BitCounter\(2)) # ((!\GenClks|BitCounter\(0)) # (!\GenClks|BitCounter[1]~DUPLICATE_q\)))) ) ) # ( !\GenClks|Equal0~0_combout\ & ( 
-- \GenClks|Add0~29_sumout\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111000011110000111100001111000011100000111100001110",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \GenClks|ALT_INV_BitCounter\(2),
	datab => \GenClks|ALT_INV_BitCounter\(0),
	datac => \GenClks|ALT_INV_Add0~29_sumout\,
	datad => \GenClks|ALT_INV_BitCounter[1]~DUPLICATE_q\,
	dataf => \GenClks|ALT_INV_Equal0~0_combout\,
	combout => \GenClks|BitCounter~1_combout\);

-- Location: FF_X15_Y64_N10
\GenClks|BitCounter[3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \GenClks|BitCounter~1_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	ena => \GenClks|ADClrc~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \GenClks|BitCounter\(3));

-- Location: MLABCELL_X15_Y64_N42
\GenClks|Add0~25\ : cyclonev_lcell_comb
-- Equation(s):
-- \GenClks|Add0~25_sumout\ = SUM(( \GenClks|BitCounter\(4) ) + ( GND ) + ( \GenClks|Add0~30\ ))
-- \GenClks|Add0~26\ = CARRY(( \GenClks|BitCounter\(4) ) + ( GND ) + ( \GenClks|Add0~30\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \GenClks|ALT_INV_BitCounter\(4),
	cin => \GenClks|Add0~30\,
	sumout => \GenClks|Add0~25_sumout\,
	cout => \GenClks|Add0~26\);

-- Location: FF_X15_Y64_N44
\GenClks|BitCounter[4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \GenClks|Add0~25_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	ena => \GenClks|ADClrc~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \GenClks|BitCounter\(4));

-- Location: MLABCELL_X15_Y64_N45
\GenClks|Add0~21\ : cyclonev_lcell_comb
-- Equation(s):
-- \GenClks|Add0~21_sumout\ = SUM(( \GenClks|BitCounter\(5) ) + ( GND ) + ( \GenClks|Add0~26\ ))
-- \GenClks|Add0~22\ = CARRY(( \GenClks|BitCounter\(5) ) + ( GND ) + ( \GenClks|Add0~26\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \GenClks|ALT_INV_BitCounter\(5),
	cin => \GenClks|Add0~26\,
	sumout => \GenClks|Add0~21_sumout\,
	cout => \GenClks|Add0~22\);

-- Location: FF_X15_Y64_N47
\GenClks|BitCounter[5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \GenClks|Add0~21_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	ena => \GenClks|ADClrc~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \GenClks|BitCounter\(5));

-- Location: MLABCELL_X15_Y64_N48
\GenClks|Add0~17\ : cyclonev_lcell_comb
-- Equation(s):
-- \GenClks|Add0~17_sumout\ = SUM(( \GenClks|BitCounter\(6) ) + ( GND ) + ( \GenClks|Add0~22\ ))
-- \GenClks|Add0~18\ = CARRY(( \GenClks|BitCounter\(6) ) + ( GND ) + ( \GenClks|Add0~22\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \GenClks|ALT_INV_BitCounter\(6),
	cin => \GenClks|Add0~22\,
	sumout => \GenClks|Add0~17_sumout\,
	cout => \GenClks|Add0~18\);

-- Location: FF_X15_Y64_N50
\GenClks|BitCounter[6]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \GenClks|Add0~17_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	ena => \GenClks|ADClrc~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \GenClks|BitCounter\(6));

-- Location: MLABCELL_X15_Y64_N51
\GenClks|Add0~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \GenClks|Add0~13_sumout\ = SUM(( \GenClks|BitCounter\(7) ) + ( GND ) + ( \GenClks|Add0~18\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \GenClks|ALT_INV_BitCounter\(7),
	cin => \GenClks|Add0~18\,
	sumout => \GenClks|Add0~13_sumout\);

-- Location: MLABCELL_X15_Y64_N6
\GenClks|BitCounter~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \GenClks|BitCounter~0_combout\ = ( \GenClks|Equal0~0_combout\ & ( (\GenClks|Add0~13_sumout\ & ((!\GenClks|BitCounter\(2)) # ((!\GenClks|BitCounter\(0)) # (!\GenClks|BitCounter\(1))))) ) ) # ( !\GenClks|Equal0~0_combout\ & ( \GenClks|Add0~13_sumout\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011111111000000001111111100000000111111100000000011111110",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \GenClks|ALT_INV_BitCounter\(2),
	datab => \GenClks|ALT_INV_BitCounter\(0),
	datac => \GenClks|ALT_INV_BitCounter\(1),
	datad => \GenClks|ALT_INV_Add0~13_sumout\,
	dataf => \GenClks|ALT_INV_Equal0~0_combout\,
	combout => \GenClks|BitCounter~0_combout\);

-- Location: FF_X15_Y64_N8
\GenClks|BitCounter[7]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \GenClks|BitCounter~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	ena => \GenClks|ADClrc~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \GenClks|BitCounter\(7));

-- Location: MLABCELL_X15_Y64_N24
\GenClks|Equal0~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \GenClks|Equal0~0_combout\ = ( !\GenClks|BitCounter\(5) & ( !\GenClks|BitCounter\(4) & ( (!\GenClks|BitCounter\(3) & (\GenClks|BitCounter\(7) & !\GenClks|BitCounter\(6))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0010000000100000000000000000000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \GenClks|ALT_INV_BitCounter\(3),
	datab => \GenClks|ALT_INV_BitCounter\(7),
	datac => \GenClks|ALT_INV_BitCounter\(6),
	datae => \GenClks|ALT_INV_BitCounter\(5),
	dataf => \GenClks|ALT_INV_BitCounter\(4),
	combout => \GenClks|Equal0~0_combout\);

-- Location: MLABCELL_X15_Y64_N18
\GenClks|ADClrc~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \GenClks|ADClrc~1_combout\ = ( \GenClks|ADClrc~q\ & ( \GenClks|BitCounter[1]~DUPLICATE_q\ & ( (!\GenClks|BitCounter\(2)) # ((!\GenClks|ADClrc~0_combout\) # ((!\GenClks|Equal0~0_combout\) # (!\GenClks|BitCounter\(0)))) ) ) ) # ( !\GenClks|ADClrc~q\ & ( 
-- \GenClks|BitCounter[1]~DUPLICATE_q\ & ( (\GenClks|BitCounter\(2) & (\GenClks|ADClrc~0_combout\ & (\GenClks|Equal0~0_combout\ & \GenClks|BitCounter\(0)))) ) ) ) # ( \GenClks|ADClrc~q\ & ( !\GenClks|BitCounter[1]~DUPLICATE_q\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000011111111111111110",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \GenClks|ALT_INV_BitCounter\(2),
	datab => \GenClks|ALT_INV_ADClrc~0_combout\,
	datac => \GenClks|ALT_INV_Equal0~0_combout\,
	datad => \GenClks|ALT_INV_BitCounter\(0),
	datae => \GenClks|ALT_INV_ADClrc~q\,
	dataf => \GenClks|ALT_INV_BitCounter[1]~DUPLICATE_q\,
	combout => \GenClks|ADClrc~1_combout\);

-- Location: FF_X15_Y64_N20
\GenClks|ADClrc\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \GenClks|ADClrc~1_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \GenClks|ADClrc~q\);

-- Location: FF_X15_Y64_N23
\TheI2sToPar|LrcDlyd\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	asdata => \GenClks|ADClrc~q\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheI2sToPar|LrcDlyd~q\);

-- Location: FF_X13_Y63_N2
\TheI2sToPar|BclkDlyd\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	asdata => \GenClks|BMclk~q\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheI2sToPar|BclkDlyd~q\);

-- Location: LABCELL_X12_Y63_N51
\TheI2sToPar|BclkRiseEdge\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheI2sToPar|BclkRiseEdge~combout\ = ( !\TheI2sToPar|BclkDlyd~q\ & ( \GenClks|BMclk~q\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011111111000000001111111100000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \GenClks|ALT_INV_BMclk~q\,
	dataf => \TheI2sToPar|ALT_INV_BclkDlyd~q\,
	combout => \TheI2sToPar|BclkRiseEdge~combout\);

-- Location: MLABCELL_X15_Y64_N54
\TheI2sToPar|State~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheI2sToPar|State~0_combout\ = ( \TheI2sToPar|BclkRiseEdge~combout\ & ( (!\TheI2sToPar|State~q\ & (!\GenClks|ADClrc~q\ $ (((!\TheI2sToPar|LrcDlyd~q\))))) # (\TheI2sToPar|State~q\ & (((!\TheI2sToPar|Equal0~1_combout\)))) ) ) # ( 
-- !\TheI2sToPar|BclkRiseEdge~combout\ & ( (!\GenClks|ADClrc~q\ $ (!\TheI2sToPar|LrcDlyd~q\)) # (\TheI2sToPar|State~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101101011111111010110101111111101011010110011000101101011001100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \GenClks|ALT_INV_ADClrc~q\,
	datab => \TheI2sToPar|ALT_INV_Equal0~1_combout\,
	datac => \TheI2sToPar|ALT_INV_LrcDlyd~q\,
	datad => \TheI2sToPar|ALT_INV_State~q\,
	dataf => \TheI2sToPar|ALT_INV_BclkRiseEdge~combout\,
	combout => \TheI2sToPar|State~0_combout\);

-- Location: FF_X15_Y64_N55
\TheI2sToPar|State\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \TheI2sToPar|State~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheI2sToPar|State~q\);

-- Location: LABCELL_X12_Y63_N0
\TheI2sToPar|NextAudioBitCtr[0]~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheI2sToPar|NextAudioBitCtr[0]~4_combout\ = ( \TheI2sToPar|BclkDlyd~q\ & ( (\TheI2sToPar|State~q\ & \TheI2sToPar|AudioBitCtr\(0)) ) ) # ( !\TheI2sToPar|BclkDlyd~q\ & ( (\TheI2sToPar|State~q\ & (!\GenClks|BMclk~q\ $ (!\TheI2sToPar|AudioBitCtr\(0)))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100001010000001010000101000000000000011110000000000001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \GenClks|ALT_INV_BMclk~q\,
	datac => \TheI2sToPar|ALT_INV_State~q\,
	datad => \TheI2sToPar|ALT_INV_AudioBitCtr\(0),
	dataf => \TheI2sToPar|ALT_INV_BclkDlyd~q\,
	combout => \TheI2sToPar|NextAudioBitCtr[0]~4_combout\);

-- Location: FF_X12_Y63_N2
\TheI2sToPar|AudioBitCtr[0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \TheI2sToPar|NextAudioBitCtr[0]~4_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheI2sToPar|AudioBitCtr\(0));

-- Location: LABCELL_X12_Y63_N45
\TheI2sToPar|NextAudioBitCtr[1]~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheI2sToPar|NextAudioBitCtr[1]~3_combout\ = ( \TheI2sToPar|BclkDlyd~q\ & ( (\TheI2sToPar|State~q\ & \TheI2sToPar|AudioBitCtr\(1)) ) ) # ( !\TheI2sToPar|BclkDlyd~q\ & ( (\TheI2sToPar|State~q\ & (!\TheI2sToPar|AudioBitCtr\(1) $ (((!\GenClks|BMclk~q\) # 
-- (\TheI2sToPar|AudioBitCtr\(0)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010000001011000001000000101100000000000011110000000000001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \GenClks|ALT_INV_BMclk~q\,
	datab => \TheI2sToPar|ALT_INV_AudioBitCtr\(0),
	datac => \TheI2sToPar|ALT_INV_State~q\,
	datad => \TheI2sToPar|ALT_INV_AudioBitCtr\(1),
	dataf => \TheI2sToPar|ALT_INV_BclkDlyd~q\,
	combout => \TheI2sToPar|NextAudioBitCtr[1]~3_combout\);

-- Location: FF_X12_Y63_N47
\TheI2sToPar|AudioBitCtr[1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \TheI2sToPar|NextAudioBitCtr[1]~3_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheI2sToPar|AudioBitCtr\(1));

-- Location: FF_X12_Y63_N46
\TheI2sToPar|AudioBitCtr[1]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \TheI2sToPar|NextAudioBitCtr[1]~3_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheI2sToPar|AudioBitCtr[1]~DUPLICATE_q\);

-- Location: FF_X12_Y63_N26
\TheI2sToPar|AudioBitCtr[2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \TheI2sToPar|NextAudioBitCtr[2]~2_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheI2sToPar|AudioBitCtr\(2));

-- Location: LABCELL_X12_Y63_N24
\TheI2sToPar|NextAudioBitCtr[2]~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheI2sToPar|NextAudioBitCtr[2]~2_combout\ = ( \TheI2sToPar|AudioBitCtr\(2) & ( \TheI2sToPar|BclkDlyd~q\ & ( \TheI2sToPar|State~q\ ) ) ) # ( \TheI2sToPar|AudioBitCtr\(2) & ( !\TheI2sToPar|BclkDlyd~q\ & ( (\TheI2sToPar|State~q\ & ((!\GenClks|BMclk~q\) # 
-- ((\TheI2sToPar|AudioBitCtr[1]~DUPLICATE_q\) # (\TheI2sToPar|AudioBitCtr\(0))))) ) ) ) # ( !\TheI2sToPar|AudioBitCtr\(2) & ( !\TheI2sToPar|BclkDlyd~q\ & ( (\GenClks|BMclk~q\ & (!\TheI2sToPar|AudioBitCtr\(0) & (\TheI2sToPar|State~q\ & 
-- !\TheI2sToPar|AudioBitCtr[1]~DUPLICATE_q\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010000000000000010110000111100000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \GenClks|ALT_INV_BMclk~q\,
	datab => \TheI2sToPar|ALT_INV_AudioBitCtr\(0),
	datac => \TheI2sToPar|ALT_INV_State~q\,
	datad => \TheI2sToPar|ALT_INV_AudioBitCtr[1]~DUPLICATE_q\,
	datae => \TheI2sToPar|ALT_INV_AudioBitCtr\(2),
	dataf => \TheI2sToPar|ALT_INV_BclkDlyd~q\,
	combout => \TheI2sToPar|NextAudioBitCtr[2]~2_combout\);

-- Location: FF_X12_Y63_N25
\TheI2sToPar|AudioBitCtr[2]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \TheI2sToPar|NextAudioBitCtr[2]~2_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheI2sToPar|AudioBitCtr[2]~DUPLICATE_q\);

-- Location: LABCELL_X12_Y63_N42
\TheI2sToPar|Equal0~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheI2sToPar|Equal0~0_combout\ = ( !\TheI2sToPar|AudioBitCtr[2]~DUPLICATE_q\ & ( (!\TheI2sToPar|AudioBitCtr\(0) & !\TheI2sToPar|AudioBitCtr\(1)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111000000000000111100000000000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheI2sToPar|ALT_INV_AudioBitCtr\(0),
	datad => \TheI2sToPar|ALT_INV_AudioBitCtr\(1),
	dataf => \TheI2sToPar|ALT_INV_AudioBitCtr[2]~DUPLICATE_q\,
	combout => \TheI2sToPar|Equal0~0_combout\);

-- Location: LABCELL_X12_Y63_N15
\TheI2sToPar|NextAudioBitCtr[3]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheI2sToPar|NextAudioBitCtr[3]~0_combout\ = ( \TheI2sToPar|BclkRiseEdge~combout\ & ( (\TheI2sToPar|State~q\ & (!\TheI2sToPar|Equal0~0_combout\ $ (!\TheI2sToPar|AudioBitCtr\(3)))) ) ) # ( !\TheI2sToPar|BclkRiseEdge~combout\ & ( (\TheI2sToPar|State~q\ & 
-- \TheI2sToPar|AudioBitCtr\(3)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001010101000000000101010100010001010001000001000101000100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheI2sToPar|ALT_INV_State~q\,
	datab => \TheI2sToPar|ALT_INV_Equal0~0_combout\,
	datad => \TheI2sToPar|ALT_INV_AudioBitCtr\(3),
	dataf => \TheI2sToPar|ALT_INV_BclkRiseEdge~combout\,
	combout => \TheI2sToPar|NextAudioBitCtr[3]~0_combout\);

-- Location: FF_X12_Y63_N16
\TheI2sToPar|AudioBitCtr[3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \TheI2sToPar|NextAudioBitCtr[3]~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheI2sToPar|AudioBitCtr\(3));

-- Location: LABCELL_X12_Y63_N12
\TheI2sToPar|NextAudioBitCtr[4]~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheI2sToPar|NextAudioBitCtr[4]~1_combout\ = ( \TheI2sToPar|AudioBitCtr\(3) & ( (!\TheI2sToPar|State~q\) # (\TheI2sToPar|AudioBitCtr\(4)) ) ) # ( !\TheI2sToPar|AudioBitCtr\(3) & ( (!\TheI2sToPar|State~q\) # (!\TheI2sToPar|AudioBitCtr\(4) $ 
-- (((!\TheI2sToPar|Equal0~0_combout\) # (!\TheI2sToPar|BclkRiseEdge~combout\)))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1010101111111110101010111111111010101010111111111010101011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheI2sToPar|ALT_INV_State~q\,
	datab => \TheI2sToPar|ALT_INV_Equal0~0_combout\,
	datac => \TheI2sToPar|ALT_INV_BclkRiseEdge~combout\,
	datad => \TheI2sToPar|ALT_INV_AudioBitCtr\(4),
	dataf => \TheI2sToPar|ALT_INV_AudioBitCtr\(3),
	combout => \TheI2sToPar|NextAudioBitCtr[4]~1_combout\);

-- Location: FF_X12_Y63_N14
\TheI2sToPar|AudioBitCtr[4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \TheI2sToPar|NextAudioBitCtr[4]~1_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheI2sToPar|AudioBitCtr\(4));

-- Location: LABCELL_X12_Y63_N48
\TheI2sToPar|Equal0~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheI2sToPar|Equal0~1_combout\ = ( !\TheI2sToPar|AudioBitCtr\(3) & ( (!\TheI2sToPar|AudioBitCtr\(0) & (!\TheI2sToPar|AudioBitCtr\(4) & (!\TheI2sToPar|AudioBitCtr\(2) & !\TheI2sToPar|AudioBitCtr\(1)))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1000000000000000100000000000000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheI2sToPar|ALT_INV_AudioBitCtr\(0),
	datab => \TheI2sToPar|ALT_INV_AudioBitCtr\(4),
	datac => \TheI2sToPar|ALT_INV_AudioBitCtr\(2),
	datad => \TheI2sToPar|ALT_INV_AudioBitCtr\(1),
	dataf => \TheI2sToPar|ALT_INV_AudioBitCtr\(3),
	combout => \TheI2sToPar|Equal0~1_combout\);

-- Location: MLABCELL_X15_Y64_N57
\TheI2sToPar|NextValL~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheI2sToPar|NextValL~0_combout\ = (!\GenClks|ADClrc~q\ & (\TheI2sToPar|Equal0~1_combout\ & (\TheI2sToPar|State~q\ & \TheI2sToPar|BclkRiseEdge~combout\)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000010000000000000001000000000000000100000000000000010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \GenClks|ALT_INV_ADClrc~q\,
	datab => \TheI2sToPar|ALT_INV_Equal0~1_combout\,
	datac => \TheI2sToPar|ALT_INV_State~q\,
	datad => \TheI2sToPar|ALT_INV_BclkRiseEdge~combout\,
	combout => \TheI2sToPar|NextValL~0_combout\);

-- Location: FF_X15_Y64_N59
\TheI2sToPar|ValL\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \TheI2sToPar|NextValL~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheI2sToPar|ValL~q\);

-- Location: LABCELL_X16_Y64_N45
\TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~0_combout\ = ( \TheI2sToPar|ValL~q\ & ( (!\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~0_combout\) # ((!\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~1_combout\) # 
-- (!\TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~q\)) ) ) # ( !\TheI2sToPar|ValL~q\ & ( (\TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~q\ & ((!\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~0_combout\) # 
-- (!\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~1_combout\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011101110000000001110111011111111111011101111111111101110",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:11:Bandpass1|ALT_INV_Equal1~0_combout\,
	datab => \TheRxFsk|Bandpasses:11:Bandpass1|ALT_INV_Equal1~1_combout\,
	datad => \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.AddressState~q\,
	dataf => \TheI2sToPar|ALT_INV_ValL~q\,
	combout => \TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~0_combout\);

-- Location: FF_X16_Y64_N47
\TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~q\);

-- Location: FF_X16_Y64_N32
\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[1]~7_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(1));

-- Location: LABCELL_X16_Y64_N42
\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[0]~8\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[0]~8_combout\ = ( \TheI2sToPar|ValL~q\ & ( (!\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(0) & ((!\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~0_combout\) # 
-- ((!\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~1_combout\) # (!\TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~q\)))) ) ) # ( !\TheI2sToPar|ValL~q\ & ( (!\TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~q\ & 
-- (((\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(0))))) # (\TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~q\ & (!\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(0) & ((!\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~0_combout\) # 
-- (!\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~1_combout\)))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111011110000000011101111000011111110000000001111111000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:11:Bandpass1|ALT_INV_Equal1~0_combout\,
	datab => \TheRxFsk|Bandpasses:11:Bandpass1|ALT_INV_Equal1~1_combout\,
	datac => \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.AddressState~q\,
	datad => \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.ReadAddressCoef\(0),
	dataf => \TheI2sToPar|ALT_INV_ValL~q\,
	combout => \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[0]~8_combout\);

-- Location: FF_X16_Y64_N44
\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[0]~8_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(0));

-- Location: LABCELL_X16_Y64_N0
\TheRxFsk|Bandpasses:0:Bandpass0|Add2~33\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:0:Bandpass0|Add2~34\ = CARRY(( \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(0) ) + ( VCC ) + ( !VCC ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000000000000011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.ReadAddressCoef\(0),
	cin => GND,
	cout => \TheRxFsk|Bandpasses:0:Bandpass0|Add2~34\);

-- Location: LABCELL_X16_Y64_N3
\TheRxFsk|Bandpasses:0:Bandpass0|Add2~29\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:0:Bandpass0|Add2~29_sumout\ = SUM(( \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(1) ) + ( GND ) + ( \TheRxFsk|Bandpasses:0:Bandpass0|Add2~34\ ))
-- \TheRxFsk|Bandpasses:0:Bandpass0|Add2~30\ = CARRY(( \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(1) ) + ( GND ) + ( \TheRxFsk|Bandpasses:0:Bandpass0|Add2~34\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.ReadAddressCoef\(1),
	cin => \TheRxFsk|Bandpasses:0:Bandpass0|Add2~34\,
	sumout => \TheRxFsk|Bandpasses:0:Bandpass0|Add2~29_sumout\,
	cout => \TheRxFsk|Bandpasses:0:Bandpass0|Add2~30\);

-- Location: LABCELL_X16_Y64_N30
\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[1]~7\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[1]~7_combout\ = ( \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(1) & ( \TheRxFsk|Bandpasses:0:Bandpass0|Add2~29_sumout\ & ( (!\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~0_combout\) # 
-- ((!\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~1_combout\) # (!\TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~q\)) ) ) ) # ( !\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(1) & ( \TheRxFsk|Bandpasses:0:Bandpass0|Add2~29_sumout\ & ( 
-- (!\TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~q\ & (((\TheI2sToPar|ValL~q\)))) # (\TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~q\ & ((!\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~0_combout\) # ((!\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~1_combout\)))) 
-- ) ) ) # ( \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(1) & ( !\TheRxFsk|Bandpasses:0:Bandpass0|Add2~29_sumout\ & ( (!\TheI2sToPar|ValL~q\ & !\TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~q\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100000000000000001111111011101111111111101110",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:11:Bandpass1|ALT_INV_Equal1~0_combout\,
	datab => \TheRxFsk|Bandpasses:11:Bandpass1|ALT_INV_Equal1~1_combout\,
	datac => \TheI2sToPar|ALT_INV_ValL~q\,
	datad => \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.AddressState~q\,
	datae => \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.ReadAddressCoef\(1),
	dataf => \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_Add2~29_sumout\,
	combout => \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[1]~7_combout\);

-- Location: FF_X16_Y64_N31
\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[1]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[1]~7_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[1]~DUPLICATE_q\);

-- Location: FF_X16_Y64_N43
\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[0]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[0]~8_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[0]~DUPLICATE_q\);

-- Location: FF_X16_Y64_N50
\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[2]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[2]~6_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[2]~DUPLICATE_q\);

-- Location: LABCELL_X16_Y64_N6
\TheRxFsk|Bandpasses:0:Bandpass0|Add2~25\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:0:Bandpass0|Add2~25_sumout\ = SUM(( \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[2]~DUPLICATE_q\ ) + ( GND ) + ( \TheRxFsk|Bandpasses:0:Bandpass0|Add2~30\ ))
-- \TheRxFsk|Bandpasses:0:Bandpass0|Add2~26\ = CARRY(( \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[2]~DUPLICATE_q\ ) + ( GND ) + ( \TheRxFsk|Bandpasses:0:Bandpass0|Add2~30\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.ReadAddressCoef[2]~DUPLICATE_q\,
	cin => \TheRxFsk|Bandpasses:0:Bandpass0|Add2~30\,
	sumout => \TheRxFsk|Bandpasses:0:Bandpass0|Add2~25_sumout\,
	cout => \TheRxFsk|Bandpasses:0:Bandpass0|Add2~26\);

-- Location: LABCELL_X16_Y64_N48
\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[2]~6\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[2]~6_combout\ = ( \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(2) & ( \TheRxFsk|Bandpasses:0:Bandpass0|Add2~25_sumout\ & ( (!\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~0_combout\) # 
-- ((!\TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~q\) # (!\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~1_combout\)) ) ) ) # ( !\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(2) & ( \TheRxFsk|Bandpasses:0:Bandpass0|Add2~25_sumout\ & ( 
-- (!\TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~q\ & (((\TheI2sToPar|ValL~q\)))) # (\TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~q\ & ((!\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~0_combout\) # ((!\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~1_combout\)))) 
-- ) ) ) # ( \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(2) & ( !\TheRxFsk|Bandpasses:0:Bandpass0|Add2~25_sumout\ & ( (!\TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~q\ & !\TheI2sToPar|ValL~q\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000110000001100000000111111001011101111111111101110",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:11:Bandpass1|ALT_INV_Equal1~0_combout\,
	datab => \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.AddressState~q\,
	datac => \TheI2sToPar|ALT_INV_ValL~q\,
	datad => \TheRxFsk|Bandpasses:11:Bandpass1|ALT_INV_Equal1~1_combout\,
	datae => \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.ReadAddressCoef\(2),
	dataf => \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_Add2~25_sumout\,
	combout => \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[2]~6_combout\);

-- Location: FF_X16_Y64_N49
\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[2]~6_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(2));

-- Location: LABCELL_X16_Y65_N30
\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:11:Bandpass1|Equal1~1_combout\ = ( !\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(2) & ( (!\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[1]~DUPLICATE_q\ & \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[0]~DUPLICATE_q\) 
-- ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011001100000000001100110000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.ReadAddressCoef[1]~DUPLICATE_q\,
	datad => \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.ReadAddressCoef[0]~DUPLICATE_q\,
	dataf => \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.ReadAddressCoef\(2),
	combout => \TheRxFsk|Bandpasses:11:Bandpass1|Equal1~1_combout\);

-- Location: FF_X16_Y64_N59
\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[6]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[6]~2_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(6));

-- Location: LABCELL_X16_Y64_N9
\TheRxFsk|Bandpasses:0:Bandpass0|Add2~21\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:0:Bandpass0|Add2~21_sumout\ = SUM(( \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(3) ) + ( GND ) + ( \TheRxFsk|Bandpasses:0:Bandpass0|Add2~26\ ))
-- \TheRxFsk|Bandpasses:0:Bandpass0|Add2~22\ = CARRY(( \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(3) ) + ( GND ) + ( \TheRxFsk|Bandpasses:0:Bandpass0|Add2~26\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.ReadAddressCoef\(3),
	cin => \TheRxFsk|Bandpasses:0:Bandpass0|Add2~26\,
	sumout => \TheRxFsk|Bandpasses:0:Bandpass0|Add2~21_sumout\,
	cout => \TheRxFsk|Bandpasses:0:Bandpass0|Add2~22\);

-- Location: LABCELL_X16_Y64_N51
\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[3]~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[3]~5_combout\ = ( \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(3) & ( \TheRxFsk|Bandpasses:0:Bandpass0|Add2~21_sumout\ & ( (!\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~0_combout\) # 
-- ((!\TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~q\) # (!\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~1_combout\)) ) ) ) # ( !\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(3) & ( \TheRxFsk|Bandpasses:0:Bandpass0|Add2~21_sumout\ & ( 
-- (!\TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~q\ & (((\TheI2sToPar|ValL~q\)))) # (\TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~q\ & ((!\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~0_combout\) # ((!\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~1_combout\)))) 
-- ) ) ) # ( \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(3) & ( !\TheRxFsk|Bandpasses:0:Bandpass0|Add2~21_sumout\ & ( (!\TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~q\ & !\TheI2sToPar|ValL~q\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000110011000000000000110010111111101111111011111110",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:11:Bandpass1|ALT_INV_Equal1~0_combout\,
	datab => \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.AddressState~q\,
	datac => \TheRxFsk|Bandpasses:11:Bandpass1|ALT_INV_Equal1~1_combout\,
	datad => \TheI2sToPar|ALT_INV_ValL~q\,
	datae => \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.ReadAddressCoef\(3),
	dataf => \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_Add2~21_sumout\,
	combout => \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[3]~5_combout\);

-- Location: FF_X16_Y64_N52
\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[3]~5_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(3));

-- Location: LABCELL_X16_Y64_N12
\TheRxFsk|Bandpasses:0:Bandpass0|Add2~17\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:0:Bandpass0|Add2~17_sumout\ = SUM(( \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(4) ) + ( GND ) + ( \TheRxFsk|Bandpasses:0:Bandpass0|Add2~22\ ))
-- \TheRxFsk|Bandpasses:0:Bandpass0|Add2~18\ = CARRY(( \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(4) ) + ( GND ) + ( \TheRxFsk|Bandpasses:0:Bandpass0|Add2~22\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.ReadAddressCoef\(4),
	cin => \TheRxFsk|Bandpasses:0:Bandpass0|Add2~22\,
	sumout => \TheRxFsk|Bandpasses:0:Bandpass0|Add2~17_sumout\,
	cout => \TheRxFsk|Bandpasses:0:Bandpass0|Add2~18\);

-- Location: LABCELL_X16_Y64_N33
\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[4]~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[4]~4_combout\ = ( \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(4) & ( \TheRxFsk|Bandpasses:0:Bandpass0|Add2~17_sumout\ & ( (!\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~0_combout\) # 
-- ((!\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~1_combout\) # (!\TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~q\)) ) ) ) # ( !\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(4) & ( \TheRxFsk|Bandpasses:0:Bandpass0|Add2~17_sumout\ & ( 
-- (!\TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~q\ & (((\TheI2sToPar|ValL~q\)))) # (\TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~q\ & ((!\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~0_combout\) # ((!\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~1_combout\)))) 
-- ) ) ) # ( \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(4) & ( !\TheRxFsk|Bandpasses:0:Bandpass0|Add2~17_sumout\ & ( (!\TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~q\ & !\TheI2sToPar|ValL~q\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100000000000000001110111111101111111011111110",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:11:Bandpass1|ALT_INV_Equal1~0_combout\,
	datab => \TheRxFsk|Bandpasses:11:Bandpass1|ALT_INV_Equal1~1_combout\,
	datac => \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.AddressState~q\,
	datad => \TheI2sToPar|ALT_INV_ValL~q\,
	datae => \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.ReadAddressCoef\(4),
	dataf => \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_Add2~17_sumout\,
	combout => \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[4]~4_combout\);

-- Location: FF_X16_Y64_N35
\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[4]~4_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(4));

-- Location: LABCELL_X16_Y64_N15
\TheRxFsk|Bandpasses:0:Bandpass0|Add2~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:0:Bandpass0|Add2~13_sumout\ = SUM(( \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(5) ) + ( GND ) + ( \TheRxFsk|Bandpasses:0:Bandpass0|Add2~18\ ))
-- \TheRxFsk|Bandpasses:0:Bandpass0|Add2~14\ = CARRY(( \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(5) ) + ( GND ) + ( \TheRxFsk|Bandpasses:0:Bandpass0|Add2~18\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.ReadAddressCoef\(5),
	cin => \TheRxFsk|Bandpasses:0:Bandpass0|Add2~18\,
	sumout => \TheRxFsk|Bandpasses:0:Bandpass0|Add2~13_sumout\,
	cout => \TheRxFsk|Bandpasses:0:Bandpass0|Add2~14\);

-- Location: LABCELL_X16_Y64_N36
\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[5]~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[5]~3_combout\ = ( \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(5) & ( \TheRxFsk|Bandpasses:0:Bandpass0|Add2~13_sumout\ & ( (!\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~0_combout\) # 
-- ((!\TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~q\) # (!\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~1_combout\)) ) ) ) # ( !\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(5) & ( \TheRxFsk|Bandpasses:0:Bandpass0|Add2~13_sumout\ & ( 
-- (!\TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~q\ & (((\TheI2sToPar|ValL~q\)))) # (\TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~q\ & ((!\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~0_combout\) # ((!\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~1_combout\)))) 
-- ) ) ) # ( \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(5) & ( !\TheRxFsk|Bandpasses:0:Bandpass0|Add2~13_sumout\ & ( (!\TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~q\ & !\TheI2sToPar|ValL~q\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000110000001100000000111111001011101111111111101110",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:11:Bandpass1|ALT_INV_Equal1~0_combout\,
	datab => \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.AddressState~q\,
	datac => \TheI2sToPar|ALT_INV_ValL~q\,
	datad => \TheRxFsk|Bandpasses:11:Bandpass1|ALT_INV_Equal1~1_combout\,
	datae => \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.ReadAddressCoef\(5),
	dataf => \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_Add2~13_sumout\,
	combout => \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[5]~3_combout\);

-- Location: FF_X16_Y64_N38
\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[5]~3_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(5));

-- Location: LABCELL_X16_Y64_N18
\TheRxFsk|Bandpasses:0:Bandpass0|Add2~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:0:Bandpass0|Add2~9_sumout\ = SUM(( \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(6) ) + ( GND ) + ( \TheRxFsk|Bandpasses:0:Bandpass0|Add2~14\ ))
-- \TheRxFsk|Bandpasses:0:Bandpass0|Add2~10\ = CARRY(( \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(6) ) + ( GND ) + ( \TheRxFsk|Bandpasses:0:Bandpass0|Add2~14\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.ReadAddressCoef\(6),
	cin => \TheRxFsk|Bandpasses:0:Bandpass0|Add2~14\,
	sumout => \TheRxFsk|Bandpasses:0:Bandpass0|Add2~9_sumout\,
	cout => \TheRxFsk|Bandpasses:0:Bandpass0|Add2~10\);

-- Location: LABCELL_X16_Y64_N57
\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[6]~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[6]~2_combout\ = ( \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(6) & ( \TheRxFsk|Bandpasses:0:Bandpass0|Add2~9_sumout\ & ( (!\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~0_combout\) # 
-- ((!\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~1_combout\) # (!\TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~q\)) ) ) ) # ( !\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(6) & ( \TheRxFsk|Bandpasses:0:Bandpass0|Add2~9_sumout\ & ( 
-- (!\TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~q\ & (((\TheI2sToPar|ValL~q\)))) # (\TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~q\ & ((!\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~0_combout\) # ((!\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~1_combout\)))) 
-- ) ) ) # ( \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(6) & ( !\TheRxFsk|Bandpasses:0:Bandpass0|Add2~9_sumout\ & ( (!\TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~q\ & !\TheI2sToPar|ValL~q\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100000000000000001110111111101111111011111110",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:11:Bandpass1|ALT_INV_Equal1~0_combout\,
	datab => \TheRxFsk|Bandpasses:11:Bandpass1|ALT_INV_Equal1~1_combout\,
	datac => \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.AddressState~q\,
	datad => \TheI2sToPar|ALT_INV_ValL~q\,
	datae => \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.ReadAddressCoef\(6),
	dataf => \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_Add2~9_sumout\,
	combout => \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[6]~2_combout\);

-- Location: FF_X16_Y64_N58
\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[6]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[6]~2_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[6]~DUPLICATE_q\);

-- Location: FF_X16_Y64_N34
\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[4]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[4]~4_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[4]~DUPLICATE_q\);

-- Location: FF_X16_Y64_N41
\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[7]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[7]~1_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(7));

-- Location: LABCELL_X16_Y64_N21
\TheRxFsk|Bandpasses:0:Bandpass0|Add2~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:0:Bandpass0|Add2~5_sumout\ = SUM(( \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(7) ) + ( GND ) + ( \TheRxFsk|Bandpasses:0:Bandpass0|Add2~10\ ))
-- \TheRxFsk|Bandpasses:0:Bandpass0|Add2~6\ = CARRY(( \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(7) ) + ( GND ) + ( \TheRxFsk|Bandpasses:0:Bandpass0|Add2~10\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.ReadAddressCoef\(7),
	cin => \TheRxFsk|Bandpasses:0:Bandpass0|Add2~10\,
	sumout => \TheRxFsk|Bandpasses:0:Bandpass0|Add2~5_sumout\,
	cout => \TheRxFsk|Bandpasses:0:Bandpass0|Add2~6\);

-- Location: LABCELL_X16_Y64_N39
\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[7]~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[7]~1_combout\ = ( \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(7) & ( \TheRxFsk|Bandpasses:0:Bandpass0|Add2~5_sumout\ & ( (!\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~0_combout\) # 
-- ((!\TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~q\) # (!\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~1_combout\)) ) ) ) # ( !\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(7) & ( \TheRxFsk|Bandpasses:0:Bandpass0|Add2~5_sumout\ & ( 
-- (!\TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~q\ & (((\TheI2sToPar|ValL~q\)))) # (\TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~q\ & ((!\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~0_combout\) # ((!\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~1_combout\)))) 
-- ) ) ) # ( \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(7) & ( !\TheRxFsk|Bandpasses:0:Bandpass0|Add2~5_sumout\ & ( (!\TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~q\ & !\TheI2sToPar|ValL~q\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000110011000000000000110010111111101111111011111110",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:11:Bandpass1|ALT_INV_Equal1~0_combout\,
	datab => \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.AddressState~q\,
	datac => \TheRxFsk|Bandpasses:11:Bandpass1|ALT_INV_Equal1~1_combout\,
	datad => \TheI2sToPar|ALT_INV_ValL~q\,
	datae => \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.ReadAddressCoef\(7),
	dataf => \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_Add2~5_sumout\,
	combout => \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[7]~1_combout\);

-- Location: FF_X16_Y64_N40
\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[7]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[7]~1_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[7]~DUPLICATE_q\);

-- Location: LABCELL_X16_Y64_N24
\TheRxFsk|Bandpasses:0:Bandpass0|Add2~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:0:Bandpass0|Add2~1_sumout\ = SUM(( \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(8) ) + ( GND ) + ( \TheRxFsk|Bandpasses:0:Bandpass0|Add2~6\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.ReadAddressCoef\(8),
	cin => \TheRxFsk|Bandpasses:0:Bandpass0|Add2~6\,
	sumout => \TheRxFsk|Bandpasses:0:Bandpass0|Add2~1_sumout\);

-- Location: LABCELL_X16_Y64_N54
\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[8]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[8]~0_combout\ = ( \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(8) & ( \TheRxFsk|Bandpasses:0:Bandpass0|Add2~1_sumout\ & ( (!\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~0_combout\) # 
-- ((!\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~1_combout\) # (!\TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~q\)) ) ) ) # ( !\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(8) & ( \TheRxFsk|Bandpasses:0:Bandpass0|Add2~1_sumout\ & ( 
-- (!\TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~q\ & (((\TheI2sToPar|ValL~q\)))) # (\TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~q\ & ((!\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~0_combout\) # ((!\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~1_combout\)))) 
-- ) ) ) # ( \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(8) & ( !\TheRxFsk|Bandpasses:0:Bandpass0|Add2~1_sumout\ & ( (!\TheI2sToPar|ValL~q\ & !\TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~q\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100000000000000001111111011101111111111101110",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:11:Bandpass1|ALT_INV_Equal1~0_combout\,
	datab => \TheRxFsk|Bandpasses:11:Bandpass1|ALT_INV_Equal1~1_combout\,
	datac => \TheI2sToPar|ALT_INV_ValL~q\,
	datad => \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.AddressState~q\,
	datae => \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.ReadAddressCoef\(8),
	dataf => \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_Add2~1_sumout\,
	combout => \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[8]~0_combout\);

-- Location: FF_X16_Y64_N55
\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[8]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[8]~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(8));

-- Location: FF_X16_Y64_N37
\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[5]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[5]~3_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[5]~DUPLICATE_q\);

-- Location: MLABCELL_X25_Y65_N27
\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:11:Bandpass1|Equal1~0_combout\ = ( !\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(3) & ( !\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[5]~DUPLICATE_q\ & ( 
-- (!\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[6]~DUPLICATE_q\ & (!\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[4]~DUPLICATE_q\ & (!\TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef[7]~DUPLICATE_q\ & 
-- \TheRxFsk|Bandpasses:0:Bandpass0|R.ReadAddressCoef\(8)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000010000000000000000000000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.ReadAddressCoef[6]~DUPLICATE_q\,
	datab => \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.ReadAddressCoef[4]~DUPLICATE_q\,
	datac => \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.ReadAddressCoef[7]~DUPLICATE_q\,
	datad => \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.ReadAddressCoef\(8),
	datae => \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.ReadAddressCoef\(3),
	dataf => \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.ReadAddressCoef[5]~DUPLICATE_q\,
	combout => \TheRxFsk|Bandpasses:11:Bandpass1|Equal1~0_combout\);

-- Location: FF_X25_Y64_N35
\TheRxFsk|Bandpasses:11:Bandpass0|R.SumState.SumValid\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	asdata => \TheRxFsk|Bandpasses:11:Bandpass0|R.SumState.SumWait2~q\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:11:Bandpass0|R.SumState.SumValid~q\);

-- Location: MLABCELL_X21_Y64_N39
\TheRxFsk|Bandpasses:11:Bandpass0|Selector0~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:11:Bandpass0|Selector0~0_combout\ = ( \TheRxFsk|Bandpasses:11:Bandpass0|R.SumState.Idle~q\ & ( \TheI2sToPar|ValL~q\ & ( !\TheRxFsk|Bandpasses:11:Bandpass0|R.SumState.SumValid~q\ ) ) ) # ( 
-- !\TheRxFsk|Bandpasses:11:Bandpass0|R.SumState.Idle~q\ & ( \TheI2sToPar|ValL~q\ & ( !\TheRxFsk|Bandpasses:11:Bandpass0|R.SumState.SumValid~q\ ) ) ) # ( \TheRxFsk|Bandpasses:11:Bandpass0|R.SumState.Idle~q\ & ( !\TheI2sToPar|ValL~q\ & ( 
-- !\TheRxFsk|Bandpasses:11:Bandpass0|R.SumState.SumValid~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000101010101010101010101010101010101010101010101010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:11:Bandpass0|ALT_INV_R.SumState.SumValid~q\,
	datae => \TheRxFsk|Bandpasses:11:Bandpass0|ALT_INV_R.SumState.Idle~q\,
	dataf => \TheI2sToPar|ALT_INV_ValL~q\,
	combout => \TheRxFsk|Bandpasses:11:Bandpass0|Selector0~0_combout\);

-- Location: FF_X21_Y64_N40
\TheRxFsk|Bandpasses:11:Bandpass0|R.SumState.Idle\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:11:Bandpass0|Selector0~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:11:Bandpass0|R.SumState.Idle~q\);

-- Location: LABCELL_X13_Y64_N9
\TheRxFsk|Bandpasses:11:Bandpass0|Selector1~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:11:Bandpass0|Selector1~0_combout\ = ( \TheI2sToPar|ValL~q\ & ( !\TheRxFsk|Bandpasses:11:Bandpass0|R.SumState.Idle~q\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011110000111100001111000011110000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:11:Bandpass0|ALT_INV_R.SumState.Idle~q\,
	dataf => \TheI2sToPar|ALT_INV_ValL~q\,
	combout => \TheRxFsk|Bandpasses:11:Bandpass0|Selector1~0_combout\);

-- Location: FF_X13_Y64_N10
\TheRxFsk|Bandpasses:11:Bandpass0|R.SumState.SumEnable\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:11:Bandpass0|Selector1~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:11:Bandpass0|R.SumState.SumEnable~q\);

-- Location: MLABCELL_X25_Y64_N57
\TheRxFsk|Bandpasses:11:Bandpass0|Selector2~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:11:Bandpass0|Selector2~0_combout\ = ( \TheRxFsk|Bandpasses:11:Bandpass1|Equal1~0_combout\ & ( ((!\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~1_combout\ & \TheRxFsk|Bandpasses:11:Bandpass0|R.SumState.SumSelect~q\)) # 
-- (\TheRxFsk|Bandpasses:11:Bandpass0|R.SumState.SumEnable~q\) ) ) # ( !\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~0_combout\ & ( (\TheRxFsk|Bandpasses:11:Bandpass0|R.SumState.SumSelect~q\) # (\TheRxFsk|Bandpasses:11:Bandpass0|R.SumState.SumEnable~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111111111111000011111111111100001111101011110000111110101111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:11:Bandpass1|ALT_INV_Equal1~1_combout\,
	datac => \TheRxFsk|Bandpasses:11:Bandpass0|ALT_INV_R.SumState.SumEnable~q\,
	datad => \TheRxFsk|Bandpasses:11:Bandpass0|ALT_INV_R.SumState.SumSelect~q\,
	dataf => \TheRxFsk|Bandpasses:11:Bandpass1|ALT_INV_Equal1~0_combout\,
	combout => \TheRxFsk|Bandpasses:11:Bandpass0|Selector2~0_combout\);

-- Location: FF_X25_Y64_N59
\TheRxFsk|Bandpasses:11:Bandpass0|R.SumState.SumSelect\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:11:Bandpass0|Selector2~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:11:Bandpass0|R.SumState.SumSelect~q\);

-- Location: MLABCELL_X25_Y64_N36
\TheRxFsk|Bandpasses:11:Bandpass0|Selector3~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:11:Bandpass0|Selector3~0_combout\ = ( \TheRxFsk|Bandpasses:11:Bandpass0|R.SumState.SumSelect~q\ & ( (\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~0_combout\ & \TheRxFsk|Bandpasses:11:Bandpass1|Equal1~1_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000011000000110000001100000011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:11:Bandpass1|ALT_INV_Equal1~0_combout\,
	datac => \TheRxFsk|Bandpasses:11:Bandpass1|ALT_INV_Equal1~1_combout\,
	dataf => \TheRxFsk|Bandpasses:11:Bandpass0|ALT_INV_R.SumState.SumSelect~q\,
	combout => \TheRxFsk|Bandpasses:11:Bandpass0|Selector3~0_combout\);

-- Location: FF_X25_Y64_N38
\TheRxFsk|Bandpasses:11:Bandpass0|R.SumState.SumWait1\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:11:Bandpass0|Selector3~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:11:Bandpass0|R.SumState.SumWait1~q\);

-- Location: FF_X25_Y64_N50
\TheRxFsk|Bandpasses:11:Bandpass0|R.SumState.SumWait2\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	asdata => \TheRxFsk|Bandpasses:11:Bandpass0|R.SumState.SumWait1~q\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:11:Bandpass0|R.SumState.SumWait2~q\);

-- Location: MLABCELL_X25_Y64_N12
\TheRxFsk|Bandpasses:11:Bandpass0|Selector8~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:11:Bandpass0|Selector8~0_combout\ = ((!\TheRxFsk|Bandpasses:11:Bandpass0|R.SumState.SumValid~q\ & \TheRxFsk|Bandpasses:11:Bandpass0|R.ValWet~q\)) # (\TheRxFsk|Bandpasses:11:Bandpass0|R.SumState.SumWait2~q\)

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010111110101010101011111010101010101111101010101010111110101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:11:Bandpass0|ALT_INV_R.SumState.SumWait2~q\,
	datac => \TheRxFsk|Bandpasses:11:Bandpass0|ALT_INV_R.SumState.SumValid~q\,
	datad => \TheRxFsk|Bandpasses:11:Bandpass0|ALT_INV_R.ValWet~q\,
	combout => \TheRxFsk|Bandpasses:11:Bandpass0|Selector8~0_combout\);

-- Location: FF_X25_Y64_N13
\TheRxFsk|Bandpasses:11:Bandpass0|R.ValWet\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:11:Bandpass0|Selector8~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:11:Bandpass0|R.ValWet~q\);

-- Location: MLABCELL_X28_Y64_N36
\TheRxFsk|Lowpass|R.AddressState~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|R.AddressState~0_combout\ = ( \TheRxFsk|Bandpasses:11:Bandpass0|R.ValWet~q\ & ( (!\TheRxFsk|Lowpass|CoefMemory~0_combout\) # ((!\TheRxFsk|Lowpass|Equal1~0_combout\) # (!\TheRxFsk|Lowpass|R.AddressState~q\)) ) ) # ( 
-- !\TheRxFsk|Bandpasses:11:Bandpass0|R.ValWet~q\ & ( (\TheRxFsk|Lowpass|R.AddressState~q\ & ((!\TheRxFsk|Lowpass|CoefMemory~0_combout\) # (!\TheRxFsk|Lowpass|Equal1~0_combout\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011101110000000001110111011111111111011101111111111101110",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_CoefMemory~0_combout\,
	datab => \TheRxFsk|Lowpass|ALT_INV_Equal1~0_combout\,
	datad => \TheRxFsk|Lowpass|ALT_INV_R.AddressState~q\,
	dataf => \TheRxFsk|Bandpasses:11:Bandpass0|ALT_INV_R.ValWet~q\,
	combout => \TheRxFsk|Lowpass|R.AddressState~0_combout\);

-- Location: FF_X28_Y64_N38
\TheRxFsk|Lowpass|R.AddressState\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|R.AddressState~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|R.AddressState~q\);

-- Location: LABCELL_X29_Y64_N30
\TheRxFsk|Lowpass|Add2~17\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add2~18\ = CARRY(( \TheRxFsk|Lowpass|R.ReadAddressCoef\(0) ) + ( VCC ) + ( !VCC ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(0),
	cin => GND,
	cout => \TheRxFsk|Lowpass|Add2~18\);

-- Location: LABCELL_X29_Y64_N33
\TheRxFsk|Lowpass|Add2~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add2~13_sumout\ = SUM(( \TheRxFsk|Lowpass|R.ReadAddressCoef\(1) ) + ( GND ) + ( \TheRxFsk|Lowpass|Add2~18\ ))
-- \TheRxFsk|Lowpass|Add2~14\ = CARRY(( \TheRxFsk|Lowpass|R.ReadAddressCoef\(1) ) + ( GND ) + ( \TheRxFsk|Lowpass|Add2~18\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(1),
	cin => \TheRxFsk|Lowpass|Add2~18\,
	sumout => \TheRxFsk|Lowpass|Add2~13_sumout\,
	cout => \TheRxFsk|Lowpass|Add2~14\);

-- Location: MLABCELL_X28_Y64_N45
\TheRxFsk|Lowpass|R.ReadAddressCoef[1]~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|R.ReadAddressCoef[1]~3_combout\ = ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & ( \TheRxFsk|Lowpass|Add2~13_sumout\ & ( (!\TheRxFsk|Lowpass|CoefMemory~0_combout\) # ((!\TheRxFsk|Lowpass|Equal1~0_combout\) # 
-- (!\TheRxFsk|Lowpass|R.AddressState~q\)) ) ) ) # ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & ( \TheRxFsk|Lowpass|Add2~13_sumout\ & ( (!\TheRxFsk|Lowpass|R.AddressState~q\ & (((\TheRxFsk|Bandpasses:11:Bandpass0|R.ValWet~q\)))) # 
-- (\TheRxFsk|Lowpass|R.AddressState~q\ & ((!\TheRxFsk|Lowpass|CoefMemory~0_combout\) # ((!\TheRxFsk|Lowpass|Equal1~0_combout\)))) ) ) ) # ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & ( !\TheRxFsk|Lowpass|Add2~13_sumout\ & ( 
-- (!\TheRxFsk|Bandpasses:11:Bandpass0|R.ValWet~q\ & !\TheRxFsk|Lowpass|R.AddressState~q\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000110011000000000000110011111110101111111111111010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_CoefMemory~0_combout\,
	datab => \TheRxFsk|Bandpasses:11:Bandpass0|ALT_INV_R.ValWet~q\,
	datac => \TheRxFsk|Lowpass|ALT_INV_Equal1~0_combout\,
	datad => \TheRxFsk|Lowpass|ALT_INV_R.AddressState~q\,
	datae => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(1),
	dataf => \TheRxFsk|Lowpass|ALT_INV_Add2~13_sumout\,
	combout => \TheRxFsk|Lowpass|R.ReadAddressCoef[1]~3_combout\);

-- Location: FF_X28_Y64_N46
\TheRxFsk|Lowpass|R.ReadAddressCoef[1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|R.ReadAddressCoef[1]~3_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|R.ReadAddressCoef\(1));

-- Location: LABCELL_X29_Y64_N36
\TheRxFsk|Lowpass|Add2~25\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add2~25_sumout\ = SUM(( \TheRxFsk|Lowpass|R.ReadAddressCoef\(2) ) + ( GND ) + ( \TheRxFsk|Lowpass|Add2~14\ ))
-- \TheRxFsk|Lowpass|Add2~26\ = CARRY(( \TheRxFsk|Lowpass|R.ReadAddressCoef\(2) ) + ( GND ) + ( \TheRxFsk|Lowpass|Add2~14\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(2),
	cin => \TheRxFsk|Lowpass|Add2~14\,
	sumout => \TheRxFsk|Lowpass|Add2~25_sumout\,
	cout => \TheRxFsk|Lowpass|Add2~26\);

-- Location: MLABCELL_X25_Y64_N51
\TheRxFsk|Lowpass|R.ReadAddressCoef[2]~6\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|R.ReadAddressCoef[2]~6_combout\ = ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & ( \TheRxFsk|Bandpasses:11:Bandpass0|R.ValWet~q\ & ( (\TheRxFsk|Lowpass|Add2~25_sumout\ & ((!\TheRxFsk|Lowpass|R.AddressState~q\) # 
-- ((!\TheRxFsk|Lowpass|CoefMemory~0_combout\) # (!\TheRxFsk|Lowpass|Equal1~0_combout\)))) ) ) ) # ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & ( \TheRxFsk|Bandpasses:11:Bandpass0|R.ValWet~q\ & ( (\TheRxFsk|Lowpass|Add2~25_sumout\ & 
-- ((!\TheRxFsk|Lowpass|R.AddressState~q\) # ((!\TheRxFsk|Lowpass|CoefMemory~0_combout\) # (!\TheRxFsk|Lowpass|Equal1~0_combout\)))) ) ) ) # ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & ( !\TheRxFsk|Bandpasses:11:Bandpass0|R.ValWet~q\ & ( 
-- (!\TheRxFsk|Lowpass|R.AddressState~q\) # ((\TheRxFsk|Lowpass|Add2~25_sumout\ & ((!\TheRxFsk|Lowpass|CoefMemory~0_combout\) # (!\TheRxFsk|Lowpass|Equal1~0_combout\)))) ) ) ) # ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & ( 
-- !\TheRxFsk|Bandpasses:11:Bandpass0|R.ValWet~q\ & ( (\TheRxFsk|Lowpass|R.AddressState~q\ & (\TheRxFsk|Lowpass|Add2~25_sumout\ & ((!\TheRxFsk|Lowpass|CoefMemory~0_combout\) # (!\TheRxFsk|Lowpass|Equal1~0_combout\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000100010000101110111011101000110011001100100011001100110010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_R.AddressState~q\,
	datab => \TheRxFsk|Lowpass|ALT_INV_Add2~25_sumout\,
	datac => \TheRxFsk|Lowpass|ALT_INV_CoefMemory~0_combout\,
	datad => \TheRxFsk|Lowpass|ALT_INV_Equal1~0_combout\,
	datae => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(2),
	dataf => \TheRxFsk|Bandpasses:11:Bandpass0|ALT_INV_R.ValWet~q\,
	combout => \TheRxFsk|Lowpass|R.ReadAddressCoef[2]~6_combout\);

-- Location: FF_X25_Y64_N52
\TheRxFsk|Lowpass|R.ReadAddressCoef[2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|R.ReadAddressCoef[2]~6_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|R.ReadAddressCoef\(2));

-- Location: LABCELL_X29_Y64_N39
\TheRxFsk|Lowpass|Add2~21\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add2~21_sumout\ = SUM(( \TheRxFsk|Lowpass|R.ReadAddressCoef\(3) ) + ( GND ) + ( \TheRxFsk|Lowpass|Add2~26\ ))
-- \TheRxFsk|Lowpass|Add2~22\ = CARRY(( \TheRxFsk|Lowpass|R.ReadAddressCoef\(3) ) + ( GND ) + ( \TheRxFsk|Lowpass|Add2~26\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(3),
	cin => \TheRxFsk|Lowpass|Add2~26\,
	sumout => \TheRxFsk|Lowpass|Add2~21_sumout\,
	cout => \TheRxFsk|Lowpass|Add2~22\);

-- Location: MLABCELL_X25_Y64_N6
\TheRxFsk|Lowpass|R.ReadAddressCoef[3]~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|R.ReadAddressCoef[3]~5_combout\ = ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & ( \TheRxFsk|Bandpasses:11:Bandpass0|R.ValWet~q\ & ( (\TheRxFsk|Lowpass|Add2~21_sumout\ & ((!\TheRxFsk|Lowpass|R.AddressState~q\) # 
-- ((!\TheRxFsk|Lowpass|CoefMemory~0_combout\) # (!\TheRxFsk|Lowpass|Equal1~0_combout\)))) ) ) ) # ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & ( \TheRxFsk|Bandpasses:11:Bandpass0|R.ValWet~q\ & ( (\TheRxFsk|Lowpass|Add2~21_sumout\ & 
-- ((!\TheRxFsk|Lowpass|R.AddressState~q\) # ((!\TheRxFsk|Lowpass|CoefMemory~0_combout\) # (!\TheRxFsk|Lowpass|Equal1~0_combout\)))) ) ) ) # ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & ( !\TheRxFsk|Bandpasses:11:Bandpass0|R.ValWet~q\ & ( 
-- (!\TheRxFsk|Lowpass|R.AddressState~q\) # ((\TheRxFsk|Lowpass|Add2~21_sumout\ & ((!\TheRxFsk|Lowpass|CoefMemory~0_combout\) # (!\TheRxFsk|Lowpass|Equal1~0_combout\)))) ) ) ) # ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & ( 
-- !\TheRxFsk|Bandpasses:11:Bandpass0|R.ValWet~q\ & ( (\TheRxFsk|Lowpass|R.AddressState~q\ & (\TheRxFsk|Lowpass|Add2~21_sumout\ & ((!\TheRxFsk|Lowpass|CoefMemory~0_combout\) # (!\TheRxFsk|Lowpass|Equal1~0_combout\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001010100101010101111111000000000111111100000000011111110",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_R.AddressState~q\,
	datab => \TheRxFsk|Lowpass|ALT_INV_CoefMemory~0_combout\,
	datac => \TheRxFsk|Lowpass|ALT_INV_Equal1~0_combout\,
	datad => \TheRxFsk|Lowpass|ALT_INV_Add2~21_sumout\,
	datae => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(3),
	dataf => \TheRxFsk|Bandpasses:11:Bandpass0|ALT_INV_R.ValWet~q\,
	combout => \TheRxFsk|Lowpass|R.ReadAddressCoef[3]~5_combout\);

-- Location: FF_X25_Y64_N7
\TheRxFsk|Lowpass|R.ReadAddressCoef[3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|R.ReadAddressCoef[3]~5_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|R.ReadAddressCoef\(3));

-- Location: LABCELL_X29_Y64_N42
\TheRxFsk|Lowpass|Add2~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add2~9_sumout\ = SUM(( \TheRxFsk|Lowpass|R.ReadAddressCoef\(4) ) + ( GND ) + ( \TheRxFsk|Lowpass|Add2~22\ ))
-- \TheRxFsk|Lowpass|Add2~10\ = CARRY(( \TheRxFsk|Lowpass|R.ReadAddressCoef\(4) ) + ( GND ) + ( \TheRxFsk|Lowpass|Add2~22\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(4),
	cin => \TheRxFsk|Lowpass|Add2~22\,
	sumout => \TheRxFsk|Lowpass|Add2~9_sumout\,
	cout => \TheRxFsk|Lowpass|Add2~10\);

-- Location: MLABCELL_X28_Y64_N42
\TheRxFsk|Lowpass|R.ReadAddressCoef[4]~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|R.ReadAddressCoef[4]~2_combout\ = ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & ( \TheRxFsk|Lowpass|Add2~9_sumout\ & ( (!\TheRxFsk|Lowpass|CoefMemory~0_combout\) # ((!\TheRxFsk|Lowpass|R.AddressState~q\) # 
-- (!\TheRxFsk|Lowpass|Equal1~0_combout\)) ) ) ) # ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & ( \TheRxFsk|Lowpass|Add2~9_sumout\ & ( (!\TheRxFsk|Lowpass|R.AddressState~q\ & (((\TheRxFsk|Bandpasses:11:Bandpass0|R.ValWet~q\)))) # 
-- (\TheRxFsk|Lowpass|R.AddressState~q\ & ((!\TheRxFsk|Lowpass|CoefMemory~0_combout\) # ((!\TheRxFsk|Lowpass|Equal1~0_combout\)))) ) ) ) # ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & ( !\TheRxFsk|Lowpass|Add2~9_sumout\ & ( 
-- (!\TheRxFsk|Bandpasses:11:Bandpass0|R.ValWet~q\ & !\TheRxFsk|Lowpass|R.AddressState~q\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000110000001100000000111111001110101111111111111010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_CoefMemory~0_combout\,
	datab => \TheRxFsk|Bandpasses:11:Bandpass0|ALT_INV_R.ValWet~q\,
	datac => \TheRxFsk|Lowpass|ALT_INV_R.AddressState~q\,
	datad => \TheRxFsk|Lowpass|ALT_INV_Equal1~0_combout\,
	datae => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(4),
	dataf => \TheRxFsk|Lowpass|ALT_INV_Add2~9_sumout\,
	combout => \TheRxFsk|Lowpass|R.ReadAddressCoef[4]~2_combout\);

-- Location: FF_X28_Y64_N44
\TheRxFsk|Lowpass|R.ReadAddressCoef[4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|R.ReadAddressCoef[4]~2_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|R.ReadAddressCoef\(4));

-- Location: LABCELL_X29_Y64_N45
\TheRxFsk|Lowpass|Add2~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add2~5_sumout\ = SUM(( \TheRxFsk|Lowpass|R.ReadAddressCoef\(5) ) + ( GND ) + ( \TheRxFsk|Lowpass|Add2~10\ ))
-- \TheRxFsk|Lowpass|Add2~6\ = CARRY(( \TheRxFsk|Lowpass|R.ReadAddressCoef\(5) ) + ( GND ) + ( \TheRxFsk|Lowpass|Add2~10\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(5),
	cin => \TheRxFsk|Lowpass|Add2~10\,
	sumout => \TheRxFsk|Lowpass|Add2~5_sumout\,
	cout => \TheRxFsk|Lowpass|Add2~6\);

-- Location: MLABCELL_X28_Y64_N51
\TheRxFsk|Lowpass|R.ReadAddressCoef[5]~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|R.ReadAddressCoef[5]~1_combout\ = ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & ( \TheRxFsk|Lowpass|Add2~5_sumout\ & ( (!\TheRxFsk|Lowpass|Equal1~0_combout\) # ((!\TheRxFsk|Lowpass|R.AddressState~q\) # 
-- (!\TheRxFsk|Lowpass|CoefMemory~0_combout\)) ) ) ) # ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & ( \TheRxFsk|Lowpass|Add2~5_sumout\ & ( (!\TheRxFsk|Lowpass|R.AddressState~q\ & (((\TheRxFsk|Bandpasses:11:Bandpass0|R.ValWet~q\)))) # 
-- (\TheRxFsk|Lowpass|R.AddressState~q\ & ((!\TheRxFsk|Lowpass|Equal1~0_combout\) # ((!\TheRxFsk|Lowpass|CoefMemory~0_combout\)))) ) ) ) # ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & ( !\TheRxFsk|Lowpass|Add2~5_sumout\ & ( 
-- (!\TheRxFsk|Bandpasses:11:Bandpass0|R.ValWet~q\ & !\TheRxFsk|Lowpass|R.AddressState~q\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000110000001100000000111111001110101111111111111010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_Equal1~0_combout\,
	datab => \TheRxFsk|Bandpasses:11:Bandpass0|ALT_INV_R.ValWet~q\,
	datac => \TheRxFsk|Lowpass|ALT_INV_R.AddressState~q\,
	datad => \TheRxFsk|Lowpass|ALT_INV_CoefMemory~0_combout\,
	datae => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(5),
	dataf => \TheRxFsk|Lowpass|ALT_INV_Add2~5_sumout\,
	combout => \TheRxFsk|Lowpass|R.ReadAddressCoef[5]~1_combout\);

-- Location: FF_X28_Y64_N52
\TheRxFsk|Lowpass|R.ReadAddressCoef[5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|R.ReadAddressCoef[5]~1_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|R.ReadAddressCoef\(5));

-- Location: MLABCELL_X28_Y65_N48
\TheRxFsk|Lowpass|CoefMemory~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|CoefMemory~0_combout\ = ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & ( (\TheRxFsk|Lowpass|R.ReadAddressCoef[6]~DUPLICATE_q\ & !\TheRxFsk|Lowpass|R.ReadAddressCoef\(4)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0100010001000100010001000100010000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef[6]~DUPLICATE_q\,
	datab => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(4),
	dataf => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(5),
	combout => \TheRxFsk|Lowpass|CoefMemory~0_combout\);

-- Location: MLABCELL_X28_Y64_N39
\TheRxFsk|Lowpass|R.ReadAddressCoef[0]~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|R.ReadAddressCoef[0]~4_combout\ = ( \TheRxFsk|Bandpasses:11:Bandpass0|R.ValWet~q\ & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & ((!\TheRxFsk|Lowpass|CoefMemory~0_combout\) # ((!\TheRxFsk|Lowpass|Equal1~0_combout\) # 
-- (!\TheRxFsk|Lowpass|R.AddressState~q\)))) ) ) # ( !\TheRxFsk|Bandpasses:11:Bandpass0|R.ValWet~q\ & ( (!\TheRxFsk|Lowpass|R.AddressState~q\ & (((\TheRxFsk|Lowpass|R.ReadAddressCoef\(0))))) # (\TheRxFsk|Lowpass|R.AddressState~q\ & 
-- (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & ((!\TheRxFsk|Lowpass|CoefMemory~0_combout\) # (!\TheRxFsk|Lowpass|Equal1~0_combout\)))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111011110000000011101111000011111110000000001111111000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_CoefMemory~0_combout\,
	datab => \TheRxFsk|Lowpass|ALT_INV_Equal1~0_combout\,
	datac => \TheRxFsk|Lowpass|ALT_INV_R.AddressState~q\,
	datad => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(0),
	dataf => \TheRxFsk|Bandpasses:11:Bandpass0|ALT_INV_R.ValWet~q\,
	combout => \TheRxFsk|Lowpass|R.ReadAddressCoef[0]~4_combout\);

-- Location: FF_X28_Y64_N40
\TheRxFsk|Lowpass|R.ReadAddressCoef[0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|R.ReadAddressCoef[0]~4_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|R.ReadAddressCoef\(0));

-- Location: LABCELL_X29_Y64_N24
\TheRxFsk|Lowpass|Equal1~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Equal1~0_combout\ = ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & (\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & !\TheRxFsk|Lowpass|R.ReadAddressCoef\(2))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000001010000000000000101000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(0),
	datac => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(1),
	datad => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(2),
	dataf => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(3),
	combout => \TheRxFsk|Lowpass|Equal1~0_combout\);

-- Location: FF_X28_Y64_N49
\TheRxFsk|Lowpass|R.ReadAddressCoef[6]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|R.ReadAddressCoef[6]~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|R.ReadAddressCoef\(6));

-- Location: LABCELL_X29_Y64_N48
\TheRxFsk|Lowpass|Add2~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add2~1_sumout\ = SUM(( \TheRxFsk|Lowpass|R.ReadAddressCoef\(6) ) + ( GND ) + ( \TheRxFsk|Lowpass|Add2~6\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(6),
	cin => \TheRxFsk|Lowpass|Add2~6\,
	sumout => \TheRxFsk|Lowpass|Add2~1_sumout\);

-- Location: MLABCELL_X28_Y64_N48
\TheRxFsk|Lowpass|R.ReadAddressCoef[6]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|R.ReadAddressCoef[6]~0_combout\ = ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(6) & ( \TheRxFsk|Lowpass|Add2~1_sumout\ & ( (!\TheRxFsk|Lowpass|Equal1~0_combout\) # ((!\TheRxFsk|Lowpass|CoefMemory~0_combout\) # 
-- (!\TheRxFsk|Lowpass|R.AddressState~q\)) ) ) ) # ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(6) & ( \TheRxFsk|Lowpass|Add2~1_sumout\ & ( (!\TheRxFsk|Lowpass|R.AddressState~q\ & (((\TheRxFsk|Bandpasses:11:Bandpass0|R.ValWet~q\)))) # 
-- (\TheRxFsk|Lowpass|R.AddressState~q\ & ((!\TheRxFsk|Lowpass|Equal1~0_combout\) # ((!\TheRxFsk|Lowpass|CoefMemory~0_combout\)))) ) ) ) # ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(6) & ( !\TheRxFsk|Lowpass|Add2~1_sumout\ & ( 
-- (!\TheRxFsk|Bandpasses:11:Bandpass0|R.ValWet~q\ & !\TheRxFsk|Lowpass|R.AddressState~q\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000110011000000000000110011111110101111111111111010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_Equal1~0_combout\,
	datab => \TheRxFsk|Bandpasses:11:Bandpass0|ALT_INV_R.ValWet~q\,
	datac => \TheRxFsk|Lowpass|ALT_INV_CoefMemory~0_combout\,
	datad => \TheRxFsk|Lowpass|ALT_INV_R.AddressState~q\,
	datae => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(6),
	dataf => \TheRxFsk|Lowpass|ALT_INV_Add2~1_sumout\,
	combout => \TheRxFsk|Lowpass|R.ReadAddressCoef[6]~0_combout\);

-- Location: FF_X28_Y64_N50
\TheRxFsk|Lowpass|R.ReadAddressCoef[6]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|R.ReadAddressCoef[6]~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|R.ReadAddressCoef[6]~DUPLICATE_q\);

-- Location: LABCELL_X29_Y65_N30
\TheRxFsk|Lowpass|CoefMemory~34\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|CoefMemory~34_combout\ = ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & (\TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & 
-- (\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & !\TheRxFsk|Lowpass|R.ReadAddressCoef\(4)))) ) ) ) # ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & 
-- ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(0) $ (\TheRxFsk|Lowpass|R.ReadAddressCoef\(1)))) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(0)) # 
-- (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(1)))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1101011000000000000000000000000000000010000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(3),
	datab => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(0),
	datac => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(1),
	datad => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(4),
	datae => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(5),
	dataf => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(2),
	combout => \TheRxFsk|Lowpass|CoefMemory~34_combout\);

-- Location: LABCELL_X29_Y65_N48
\TheRxFsk|Lowpass|CoefMemory~33\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|CoefMemory~33_combout\ = ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(4)) # 
-- ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & !\TheRxFsk|Lowpass|R.ReadAddressCoef\(3))))) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(0) $ ((\TheRxFsk|Lowpass|R.ReadAddressCoef\(3))))) ) ) ) # ( 
-- !\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & (\TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3)) # 
-- (\TheRxFsk|Lowpass|R.ReadAddressCoef\(1))))) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) $ (((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3)) # (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(4)))))) ) ) ) # ( 
-- \TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & (\TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3)) # 
-- (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(4))))) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & (\TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3)) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(0))))) ) ) ) # ( 
-- !\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) $ (\TheRxFsk|Lowpass|R.ReadAddressCoef\(4))))) # 
-- (\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(4)) # ((\TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & \TheRxFsk|Lowpass|R.ReadAddressCoef\(3))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111010100001011001000100111000100010001110101101110101111000001",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(1),
	datab => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(0),
	datac => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(3),
	datad => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(4),
	datae => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(5),
	dataf => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(2),
	combout => \TheRxFsk|Lowpass|CoefMemory~33_combout\);

-- Location: LABCELL_X29_Y65_N21
\TheRxFsk|Lowpass|CoefMemory~35\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|CoefMemory~35_combout\ = ( \TheRxFsk|Lowpass|CoefMemory~33_combout\ & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef[6]~DUPLICATE_q\) # (\TheRxFsk|Lowpass|CoefMemory~34_combout\) ) ) # ( !\TheRxFsk|Lowpass|CoefMemory~33_combout\ & ( 
-- (\TheRxFsk|Lowpass|R.ReadAddressCoef[6]~DUPLICATE_q\ & \TheRxFsk|Lowpass|CoefMemory~34_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100000101000001010000010110101111101011111010111110101111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef[6]~DUPLICATE_q\,
	datac => \TheRxFsk|Lowpass|ALT_INV_CoefMemory~34_combout\,
	dataf => \TheRxFsk|Lowpass|ALT_INV_CoefMemory~33_combout\,
	combout => \TheRxFsk|Lowpass|CoefMemory~35_combout\);

-- Location: LABCELL_X29_Y65_N12
\TheRxFsk|Lowpass|CoefMemory~31\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|CoefMemory~31_combout\ = ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & ( (\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & 
-- (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & !\TheRxFsk|Lowpass|R.ReadAddressCoef\(4)))) ) ) ) # ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & 
-- ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3)))) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & \TheRxFsk|Lowpass|R.ReadAddressCoef\(3))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1010010000000000000000000000000001000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(1),
	datab => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(0),
	datac => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(3),
	datad => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(4),
	datae => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(5),
	dataf => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(2),
	combout => \TheRxFsk|Lowpass|CoefMemory~31_combout\);

-- Location: LABCELL_X29_Y65_N6
\TheRxFsk|Lowpass|CoefMemory~30\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|CoefMemory~30_combout\ = ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & 
-- ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3)))) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(1))))) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & 
-- (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & \TheRxFsk|Lowpass|R.ReadAddressCoef\(4))) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & (\TheRxFsk|Lowpass|R.ReadAddressCoef\(3))))) ) ) ) # ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & ( 
-- \TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(4) $ (((\TheRxFsk|Lowpass|R.ReadAddressCoef\(0)) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(1)))))) # 
-- (\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & (\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & !\TheRxFsk|Lowpass|R.ReadAddressCoef\(4)))) ) ) ) # ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & ( 
-- !\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) $ (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3))))) # 
-- (\TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) $ (((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & \TheRxFsk|Lowpass|R.ReadAddressCoef\(4)))))) ) ) ) # ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & ( 
-- !\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) $ (\TheRxFsk|Lowpass|R.ReadAddressCoef\(3))))) # 
-- (\TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) $ (((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(4)) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(1)))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1000011100100001011010100001001010000100011100001100000110101001",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(1),
	datab => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(0),
	datac => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(3),
	datad => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(4),
	datae => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(5),
	dataf => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(2),
	combout => \TheRxFsk|Lowpass|CoefMemory~30_combout\);

-- Location: LABCELL_X29_Y65_N18
\TheRxFsk|Lowpass|CoefMemory~32\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|CoefMemory~32_combout\ = ( \TheRxFsk|Lowpass|CoefMemory~30_combout\ & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef[6]~DUPLICATE_q\) # (\TheRxFsk|Lowpass|CoefMemory~31_combout\) ) ) # ( !\TheRxFsk|Lowpass|CoefMemory~30_combout\ & ( 
-- (\TheRxFsk|Lowpass|R.ReadAddressCoef[6]~DUPLICATE_q\ & \TheRxFsk|Lowpass|CoefMemory~31_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000100010001000100010001000110111011101110111011101110111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef[6]~DUPLICATE_q\,
	datab => \TheRxFsk|Lowpass|ALT_INV_CoefMemory~31_combout\,
	dataf => \TheRxFsk|Lowpass|ALT_INV_CoefMemory~30_combout\,
	combout => \TheRxFsk|Lowpass|CoefMemory~32_combout\);

-- Location: LABCELL_X29_Y65_N0
\TheRxFsk|Lowpass|CoefMemory~28\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|CoefMemory~28_combout\ = ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & 
-- ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(0)) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(1))))) ) ) ) # ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & 
-- (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(0)) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(3))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1000101000000000000000000000000011010000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(1),
	datab => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(0),
	datac => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(3),
	datad => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(4),
	datae => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(5),
	dataf => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(2),
	combout => \TheRxFsk|Lowpass|CoefMemory~28_combout\);

-- Location: LABCELL_X29_Y65_N42
\TheRxFsk|Lowpass|CoefMemory~27\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|CoefMemory~27_combout\ = ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) $ 
-- (((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(0)) # (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(4)))))) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & 
-- \TheRxFsk|Lowpass|R.ReadAddressCoef\(4))) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(4)))))) ) ) ) # ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & ( 
-- (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & \TheRxFsk|Lowpass|R.ReadAddressCoef\(4))) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & 
-- (\TheRxFsk|Lowpass|R.ReadAddressCoef\(3))))) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3)))) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & 
-- (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(1))))) ) ) ) # ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) $ 
-- (((\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & !\TheRxFsk|Lowpass|R.ReadAddressCoef\(4)))))) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(4)))) # 
-- (\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(1))))) ) ) ) # ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & 
-- (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(0)) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(3))))) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) $ 
-- (((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(0)) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(1)))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1000101000101101101101101100001000110100101001100001101101101000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(1),
	datab => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(0),
	datac => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(3),
	datad => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(4),
	datae => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(5),
	dataf => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(2),
	combout => \TheRxFsk|Lowpass|CoefMemory~27_combout\);

-- Location: LABCELL_X29_Y65_N39
\TheRxFsk|Lowpass|CoefMemory~29\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|CoefMemory~29_combout\ = ( \TheRxFsk|Lowpass|CoefMemory~27_combout\ & ( (\TheRxFsk|Lowpass|R.ReadAddressCoef[6]~DUPLICATE_q\ & \TheRxFsk|Lowpass|CoefMemory~28_combout\) ) ) # ( !\TheRxFsk|Lowpass|CoefMemory~27_combout\ & ( 
-- (!\TheRxFsk|Lowpass|R.ReadAddressCoef[6]~DUPLICATE_q\) # (\TheRxFsk|Lowpass|CoefMemory~28_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1010101011111111101010101111111100000000010101010000000001010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef[6]~DUPLICATE_q\,
	datad => \TheRxFsk|Lowpass|ALT_INV_CoefMemory~28_combout\,
	dataf => \TheRxFsk|Lowpass|ALT_INV_CoefMemory~27_combout\,
	combout => \TheRxFsk|Lowpass|CoefMemory~29_combout\);

-- Location: LABCELL_X17_Y64_N24
\TheRxFsk|Lowpass|CoefMemory~25\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|CoefMemory~25_combout\ = ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & ( (\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & 
-- (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & !\TheRxFsk|Lowpass|R.ReadAddressCoef\(3)))) ) ) ) # ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & 
-- (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(1)) # (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3))))) ) ) ) # ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & ( 
-- (\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & !\TheRxFsk|Lowpass|R.ReadAddressCoef\(3)))) ) ) ) # ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & ( 
-- !\TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & \TheRxFsk|Lowpass|R.ReadAddressCoef\(3))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011000000010000000000000011000000100000000100000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(1),
	datab => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(5),
	datac => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(4),
	datad => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(3),
	datae => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(2),
	dataf => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(0),
	combout => \TheRxFsk|Lowpass|CoefMemory~25_combout\);

-- Location: LABCELL_X17_Y64_N6
\TheRxFsk|Lowpass|CoefMemory~24\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|CoefMemory~24_combout\ = ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & 
-- (\TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & \TheRxFsk|Lowpass|R.ReadAddressCoef\(3))) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3)))))) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & 
-- (((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & \TheRxFsk|Lowpass|R.ReadAddressCoef\(3))))) ) ) ) # ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & 
-- (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(1)) # (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3))))) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) $ 
-- (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) $ (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3))))) ) ) ) # ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & 
-- (((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(4))))) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & (\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & !\TheRxFsk|Lowpass|R.ReadAddressCoef\(3))) # 
-- (\TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & ((\TheRxFsk|Lowpass|R.ReadAddressCoef\(3)))))) ) ) ) # ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & 
-- ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(5)) # (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) $ (\TheRxFsk|Lowpass|R.ReadAddressCoef\(4))))) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & 
-- ((\TheRxFsk|Lowpass|R.ReadAddressCoef\(4)))) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & (\TheRxFsk|Lowpass|R.ReadAddressCoef\(5))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1110110100011011101100001010010111001001100001100100010000111000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(1),
	datab => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(5),
	datac => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(4),
	datad => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(3),
	datae => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(2),
	dataf => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(0),
	combout => \TheRxFsk|Lowpass|CoefMemory~24_combout\);

-- Location: LABCELL_X17_Y64_N18
\TheRxFsk|Lowpass|CoefMemory~26\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|CoefMemory~26_combout\ = ( \TheRxFsk|Lowpass|R.ReadAddressCoef[6]~DUPLICATE_q\ & ( \TheRxFsk|Lowpass|CoefMemory~24_combout\ & ( \TheRxFsk|Lowpass|CoefMemory~25_combout\ ) ) ) # ( !\TheRxFsk|Lowpass|R.ReadAddressCoef[6]~DUPLICATE_q\ & ( 
-- \TheRxFsk|Lowpass|CoefMemory~24_combout\ ) ) # ( \TheRxFsk|Lowpass|R.ReadAddressCoef[6]~DUPLICATE_q\ & ( !\TheRxFsk|Lowpass|CoefMemory~24_combout\ & ( \TheRxFsk|Lowpass|CoefMemory~25_combout\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000011110000111111111111111111110000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Lowpass|ALT_INV_CoefMemory~25_combout\,
	datae => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef[6]~DUPLICATE_q\,
	dataf => \TheRxFsk|Lowpass|ALT_INV_CoefMemory~24_combout\,
	combout => \TheRxFsk|Lowpass|CoefMemory~26_combout\);

-- Location: MLABCELL_X28_Y65_N0
\TheRxFsk|Lowpass|CoefMemory~21\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|CoefMemory~21_combout\ = ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & 
-- (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) $ (\TheRxFsk|Lowpass|R.ReadAddressCoef\(5))))) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & (\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) $ 
-- (\TheRxFsk|Lowpass|R.ReadAddressCoef\(5))))) ) ) ) # ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) $ 
-- (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(5)))) ) ) ) # ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & (((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(5))))) # 
-- (\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & (\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) $ (\TheRxFsk|Lowpass|R.ReadAddressCoef\(3))))) ) ) ) # ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & ( 
-- !\TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3)) # (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(5)))) # 
-- (\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & !\TheRxFsk|Lowpass|R.ReadAddressCoef\(5))))) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & 
-- (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) $ (\TheRxFsk|Lowpass|R.ReadAddressCoef\(5))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1110100010000100110011000010000100001100110000001000010000001001",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(1),
	datab => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(2),
	datac => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(3),
	datad => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(5),
	datae => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(0),
	dataf => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(4),
	combout => \TheRxFsk|Lowpass|CoefMemory~21_combout\);

-- Location: MLABCELL_X28_Y65_N42
\TheRxFsk|Lowpass|CoefMemory~22\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|CoefMemory~22_combout\ = ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & 
-- (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(2))) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & (\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & !\TheRxFsk|Lowpass|R.ReadAddressCoef\(3))))) ) ) ) # ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & ( 
-- !\TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & (\TheRxFsk|Lowpass|R.ReadAddressCoef\(1))) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & 
-- ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(2)))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101110000000000100110000000000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(1),
	datab => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(2),
	datac => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(3),
	datad => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(5),
	datae => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(0),
	dataf => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(4),
	combout => \TheRxFsk|Lowpass|CoefMemory~22_combout\);

-- Location: MLABCELL_X28_Y65_N30
\TheRxFsk|Lowpass|CoefMemory~23\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|CoefMemory~23_combout\ = ( \TheRxFsk|Lowpass|CoefMemory~22_combout\ & ( (\TheRxFsk|Lowpass|CoefMemory~21_combout\) # (\TheRxFsk|Lowpass|R.ReadAddressCoef[6]~DUPLICATE_q\) ) ) # ( !\TheRxFsk|Lowpass|CoefMemory~22_combout\ & ( 
-- (!\TheRxFsk|Lowpass|R.ReadAddressCoef[6]~DUPLICATE_q\ & \TheRxFsk|Lowpass|CoefMemory~21_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000101000001010000010100000101001011111010111110101111101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef[6]~DUPLICATE_q\,
	datac => \TheRxFsk|Lowpass|ALT_INV_CoefMemory~21_combout\,
	dataf => \TheRxFsk|Lowpass|ALT_INV_CoefMemory~22_combout\,
	combout => \TheRxFsk|Lowpass|CoefMemory~23_combout\);

-- Location: MLABCELL_X28_Y65_N12
\TheRxFsk|Lowpass|CoefMemory~18\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|CoefMemory~18_combout\ = ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & 
-- (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & \TheRxFsk|Lowpass|R.ReadAddressCoef\(5))) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(5)))))) ) ) ) # ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & ( 
-- \TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) $ ((\TheRxFsk|Lowpass|R.ReadAddressCoef\(3))))) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & 
-- (((\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & \TheRxFsk|Lowpass|R.ReadAddressCoef\(5))))) ) ) ) # ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & 
-- ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & ((\TheRxFsk|Lowpass|R.ReadAddressCoef\(5)))) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(1))))) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & 
-- ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3)) # ((\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & \TheRxFsk|Lowpass|R.ReadAddressCoef\(5))))) ) ) ) # ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & ( 
-- (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) $ (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(5))))) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) $ 
-- (((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3)) # (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(5)))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001101110110100001110001111100110000100100001110000110010000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(1),
	datab => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(2),
	datac => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(3),
	datad => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(5),
	datae => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(0),
	dataf => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(4),
	combout => \TheRxFsk|Lowpass|CoefMemory~18_combout\);

-- Location: MLABCELL_X28_Y65_N54
\TheRxFsk|Lowpass|CoefMemory~19\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|CoefMemory~19_combout\ = ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & 
-- (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & \TheRxFsk|Lowpass|R.ReadAddressCoef\(3))) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & (\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & !\TheRxFsk|Lowpass|R.ReadAddressCoef\(3))))) ) ) ) # ( 
-- !\TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) $ (((\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & 
-- !\TheRxFsk|Lowpass|R.ReadAddressCoef\(3)))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1001110000000000000110000000000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(1),
	datab => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(2),
	datac => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(3),
	datad => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(5),
	datae => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(0),
	dataf => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(4),
	combout => \TheRxFsk|Lowpass|CoefMemory~19_combout\);

-- Location: MLABCELL_X28_Y65_N51
\TheRxFsk|Lowpass|CoefMemory~20\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|CoefMemory~20_combout\ = (!\TheRxFsk|Lowpass|R.ReadAddressCoef[6]~DUPLICATE_q\ & (!\TheRxFsk|Lowpass|CoefMemory~18_combout\)) # (\TheRxFsk|Lowpass|R.ReadAddressCoef[6]~DUPLICATE_q\ & ((\TheRxFsk|Lowpass|CoefMemory~19_combout\)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1010000011110101101000001111010110100000111101011010000011110101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef[6]~DUPLICATE_q\,
	datac => \TheRxFsk|Lowpass|ALT_INV_CoefMemory~18_combout\,
	datad => \TheRxFsk|Lowpass|ALT_INV_CoefMemory~19_combout\,
	combout => \TheRxFsk|Lowpass|CoefMemory~20_combout\);

-- Location: LABCELL_X29_Y65_N54
\TheRxFsk|Lowpass|CoefMemory~16\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|CoefMemory~16_combout\ = ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & ( (\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & 
-- !\TheRxFsk|Lowpass|R.ReadAddressCoef\(4))) ) ) ) # ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & ( (\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & 
-- ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(1)) # (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(0))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111000000000000000000000000001010000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(1),
	datab => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(0),
	datac => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(3),
	datad => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(4),
	datae => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(5),
	dataf => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(2),
	combout => \TheRxFsk|Lowpass|CoefMemory~16_combout\);

-- Location: LABCELL_X29_Y65_N24
\TheRxFsk|Lowpass|CoefMemory~15\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|CoefMemory~15_combout\ = ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & (((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(4)) # 
-- (\TheRxFsk|Lowpass|R.ReadAddressCoef\(0))))) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(0) $ (((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & \TheRxFsk|Lowpass|R.ReadAddressCoef\(4)))))) ) ) ) # ( 
-- !\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(0)) # 
-- (\TheRxFsk|Lowpass|R.ReadAddressCoef\(3))))) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(0) $ (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3))))) ) ) ) # ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & ( 
-- !\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3))) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & 
-- (\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & \TheRxFsk|Lowpass|R.ReadAddressCoef\(4))))) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(0) $ ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3))))) ) ) ) # ( 
-- !\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) $ (((\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & 
-- \TheRxFsk|Lowpass|R.ReadAddressCoef\(4))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111000010110100100101001001011010001010001111001111110000110110",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(1),
	datab => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(0),
	datac => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(3),
	datad => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(4),
	datae => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(5),
	dataf => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(2),
	combout => \TheRxFsk|Lowpass|CoefMemory~15_combout\);

-- Location: LABCELL_X29_Y65_N36
\TheRxFsk|Lowpass|CoefMemory~17\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|CoefMemory~17_combout\ = ( \TheRxFsk|Lowpass|CoefMemory~15_combout\ & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef[6]~DUPLICATE_q\) # (\TheRxFsk|Lowpass|CoefMemory~16_combout\) ) ) # ( !\TheRxFsk|Lowpass|CoefMemory~15_combout\ & ( 
-- (\TheRxFsk|Lowpass|R.ReadAddressCoef[6]~DUPLICATE_q\ & \TheRxFsk|Lowpass|CoefMemory~16_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100000101000001010000010110101111101011111010111110101111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef[6]~DUPLICATE_q\,
	datac => \TheRxFsk|Lowpass|ALT_INV_CoefMemory~16_combout\,
	dataf => \TheRxFsk|Lowpass|ALT_INV_CoefMemory~15_combout\,
	combout => \TheRxFsk|Lowpass|CoefMemory~17_combout\);

-- Location: LABCELL_X29_Y64_N3
\TheRxFsk|Lowpass|CoefMemory~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|CoefMemory~13_combout\ = ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & (((\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & 
-- \TheRxFsk|Lowpass|R.ReadAddressCoef\(1))))) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(0)) # (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(1))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011000000101100000000000000000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(0),
	datab => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(3),
	datac => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(2),
	datad => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(1),
	datae => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(4),
	dataf => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(5),
	combout => \TheRxFsk|Lowpass|CoefMemory~13_combout\);

-- Location: LABCELL_X29_Y64_N18
\TheRxFsk|Lowpass|CoefMemory~12\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|CoefMemory~12_combout\ = ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & (((\TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & 
-- \TheRxFsk|Lowpass|R.ReadAddressCoef\(3))))) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(0)))) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & 
-- (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(2))))) ) ) ) # ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) $ (((\TheRxFsk|Lowpass|R.ReadAddressCoef\(2)) # 
-- (\TheRxFsk|Lowpass|R.ReadAddressCoef\(5)))) ) ) ) # ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(5)) # 
-- ((\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & \TheRxFsk|Lowpass|R.ReadAddressCoef\(3))))) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) $ (((\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & 
-- !\TheRxFsk|Lowpass|R.ReadAddressCoef\(2)))))) ) ) ) # ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & 
-- ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(2)) # (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(0)))) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & !\TheRxFsk|Lowpass|R.ReadAddressCoef\(0))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1110100000000000101010111011010010001000011101110101000001001110",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(5),
	datab => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(2),
	datac => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(0),
	datad => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(3),
	datae => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(4),
	dataf => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(1),
	combout => \TheRxFsk|Lowpass|CoefMemory~12_combout\);

-- Location: LABCELL_X29_Y64_N15
\TheRxFsk|Lowpass|CoefMemory~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|CoefMemory~14_combout\ = ( \TheRxFsk|Lowpass|CoefMemory~12_combout\ & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(6)) # (\TheRxFsk|Lowpass|CoefMemory~13_combout\) ) ) # ( !\TheRxFsk|Lowpass|CoefMemory~12_combout\ & ( 
-- (\TheRxFsk|Lowpass|CoefMemory~13_combout\ & \TheRxFsk|Lowpass|R.ReadAddressCoef\(6)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001010101000000000101010111111111010101011111111101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_CoefMemory~13_combout\,
	datad => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(6),
	dataf => \TheRxFsk|Lowpass|ALT_INV_CoefMemory~12_combout\,
	combout => \TheRxFsk|Lowpass|CoefMemory~14_combout\);

-- Location: LABCELL_X29_Y64_N6
\TheRxFsk|Lowpass|CoefMemory~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|CoefMemory~9_combout\ = ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(2))) # 
-- (\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & (\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & !\TheRxFsk|Lowpass|R.ReadAddressCoef\(3))) ) ) ) # ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & ( 
-- (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3)))) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & (\TheRxFsk|Lowpass|R.ReadAddressCoef\(5))) ) ) ) # ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & ( 
-- !\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) $ ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(2))))) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & 
-- (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) $ (((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & !\TheRxFsk|Lowpass|R.ReadAddressCoef\(2)))))) ) ) ) # ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & ( 
-- (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(2)) # (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(0))))) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & 
-- ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & ((\TheRxFsk|Lowpass|R.ReadAddressCoef\(3)) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(0)))) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3)))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1011110101000100011001110110100011011101000100011001100110001000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(5),
	datab => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(2),
	datac => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(0),
	datad => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(3),
	datae => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(4),
	dataf => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(1),
	combout => \TheRxFsk|Lowpass|CoefMemory~9_combout\);

-- Location: LABCELL_X29_Y64_N0
\TheRxFsk|Lowpass|CoefMemory~10\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|CoefMemory~10_combout\ = ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & (((\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & 
-- \TheRxFsk|Lowpass|R.ReadAddressCoef\(2))))) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(0)) # (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(1))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001000001100000000000000000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(0),
	datab => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(3),
	datac => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(1),
	datad => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(2),
	datae => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(4),
	dataf => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(5),
	combout => \TheRxFsk|Lowpass|CoefMemory~10_combout\);

-- Location: LABCELL_X29_Y64_N54
\TheRxFsk|Lowpass|CoefMemory~11\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|CoefMemory~11_combout\ = (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(6) & (\TheRxFsk|Lowpass|CoefMemory~9_combout\)) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(6) & ((\TheRxFsk|Lowpass|CoefMemory~10_combout\)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001100001111001100110000111100110011000011110011001100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Lowpass|ALT_INV_CoefMemory~9_combout\,
	datac => \TheRxFsk|Lowpass|ALT_INV_CoefMemory~10_combout\,
	datad => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(6),
	combout => \TheRxFsk|Lowpass|CoefMemory~11_combout\);

-- Location: MLABCELL_X28_Y65_N36
\TheRxFsk|Lowpass|CoefMemory~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|CoefMemory~2_combout\ = ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) $ 
-- (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(5))))) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & (\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & !\TheRxFsk|Lowpass|R.ReadAddressCoef\(5)))) ) ) ) # ( 
-- !\TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) $ (((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(1)) # 
-- (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(2)))))) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(1)) # (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(2))))) ) ) ) # ( 
-- \TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & (((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & !\TheRxFsk|Lowpass|R.ReadAddressCoef\(5))))) # 
-- (\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & (\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & (\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & \TheRxFsk|Lowpass|R.ReadAddressCoef\(5)))) ) ) ) # ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & ( 
-- !\TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(1)) # (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(2))))) # 
-- (\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & (\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & (\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & \TheRxFsk|Lowpass|R.ReadAddressCoef\(5)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1110000000000001110000000000000100011110111000000001110011000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(1),
	datab => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(2),
	datac => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(3),
	datad => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(5),
	datae => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(0),
	dataf => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(4),
	combout => \TheRxFsk|Lowpass|CoefMemory~2_combout\);

-- Location: MLABCELL_X28_Y65_N18
\TheRxFsk|Lowpass|CoefMemory~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|CoefMemory~1_combout\ = (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & (\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(1)) # (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(0))))) # 
-- (\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & (\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3)))))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000111001000000100011100100000010001110010000001000111001000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(1),
	datab => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(2),
	datac => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(0),
	datad => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(3),
	combout => \TheRxFsk|Lowpass|CoefMemory~1_combout\);

-- Location: MLABCELL_X28_Y65_N33
\TheRxFsk|Lowpass|CoefMemory~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|CoefMemory~3_combout\ = ( \TheRxFsk|Lowpass|CoefMemory~1_combout\ & ( ((!\TheRxFsk|Lowpass|R.ReadAddressCoef[6]~DUPLICATE_q\ & \TheRxFsk|Lowpass|CoefMemory~2_combout\)) # (\TheRxFsk|Lowpass|CoefMemory~0_combout\) ) ) # ( 
-- !\TheRxFsk|Lowpass|CoefMemory~1_combout\ & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef[6]~DUPLICATE_q\ & \TheRxFsk|Lowpass|CoefMemory~2_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000010101010000000001010101000001111101011110000111110101111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef[6]~DUPLICATE_q\,
	datac => \TheRxFsk|Lowpass|ALT_INV_CoefMemory~0_combout\,
	datad => \TheRxFsk|Lowpass|ALT_INV_CoefMemory~2_combout\,
	dataf => \TheRxFsk|Lowpass|ALT_INV_CoefMemory~1_combout\,
	combout => \TheRxFsk|Lowpass|CoefMemory~3_combout\);

-- Location: MLABCELL_X28_Y65_N21
\TheRxFsk|Lowpass|CoefMemory~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|CoefMemory~4_combout\ = (\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & (\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & ((\TheRxFsk|Lowpass|R.ReadAddressCoef\(0)) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(1)))))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000010011000000000001001100000000000100110000000000010011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(1),
	datab => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(2),
	datac => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(0),
	datad => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(3),
	combout => \TheRxFsk|Lowpass|CoefMemory~4_combout\);

-- Location: MLABCELL_X28_Y65_N24
\TheRxFsk|Lowpass|CoefMemory~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|CoefMemory~5_combout\ = ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & ( (\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & (\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & \TheRxFsk|Lowpass|R.ReadAddressCoef\(1))) ) ) # ( 
-- !\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & ( ((\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & ((\TheRxFsk|Lowpass|R.ReadAddressCoef\(0)) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(1))))) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(3)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101011101110111010101110111011100000001000000010000000100000001",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(3),
	datab => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(2),
	datac => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(1),
	datad => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(0),
	dataf => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(5),
	combout => \TheRxFsk|Lowpass|CoefMemory~5_combout\);

-- Location: MLABCELL_X28_Y65_N6
\TheRxFsk|Lowpass|CoefMemory~6\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|CoefMemory~6_combout\ = ( \TheRxFsk|Lowpass|CoefMemory~4_combout\ & ( \TheRxFsk|Lowpass|CoefMemory~5_combout\ & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef[6]~DUPLICATE_q\ & 
-- ((\TheRxFsk|Lowpass|R.ReadAddressCoef\(4)))) # (\TheRxFsk|Lowpass|R.ReadAddressCoef[6]~DUPLICATE_q\ & (\TheRxFsk|Lowpass|CoefMemory~1_combout\ & !\TheRxFsk|Lowpass|R.ReadAddressCoef\(4))))) ) ) ) # ( !\TheRxFsk|Lowpass|CoefMemory~4_combout\ & ( 
-- \TheRxFsk|Lowpass|CoefMemory~5_combout\ & ( (\TheRxFsk|Lowpass|R.ReadAddressCoef[6]~DUPLICATE_q\ & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & (\TheRxFsk|Lowpass|CoefMemory~1_combout\ & !\TheRxFsk|Lowpass|R.ReadAddressCoef\(4)))) ) ) ) # ( 
-- \TheRxFsk|Lowpass|CoefMemory~4_combout\ & ( !\TheRxFsk|Lowpass|CoefMemory~5_combout\ & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef[6]~DUPLICATE_q\ & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(5)) # ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(4))))) # 
-- (\TheRxFsk|Lowpass|R.ReadAddressCoef[6]~DUPLICATE_q\ & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & (\TheRxFsk|Lowpass|CoefMemory~1_combout\ & !\TheRxFsk|Lowpass|R.ReadAddressCoef\(4)))) ) ) ) # ( !\TheRxFsk|Lowpass|CoefMemory~4_combout\ & ( 
-- !\TheRxFsk|Lowpass|CoefMemory~5_combout\ & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef[6]~DUPLICATE_q\) # ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) & \TheRxFsk|Lowpass|CoefMemory~1_combout\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1010111000000000101011101000100000000100000000000000010010001000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef[6]~DUPLICATE_q\,
	datab => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(5),
	datac => \TheRxFsk|Lowpass|ALT_INV_CoefMemory~1_combout\,
	datad => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(4),
	datae => \TheRxFsk|Lowpass|ALT_INV_CoefMemory~4_combout\,
	dataf => \TheRxFsk|Lowpass|ALT_INV_CoefMemory~5_combout\,
	combout => \TheRxFsk|Lowpass|CoefMemory~6_combout\);

-- Location: MLABCELL_X28_Y65_N27
\TheRxFsk|Lowpass|CoefMemory~7\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|CoefMemory~7_combout\ = ( \TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & ( (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) $ (((\TheRxFsk|Lowpass|R.ReadAddressCoef[6]~DUPLICATE_q\))))) # 
-- (\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(0) & \TheRxFsk|Lowpass|R.ReadAddressCoef[6]~DUPLICATE_q\))) ) ) # ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(1) & ( 
-- (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & (!\TheRxFsk|Lowpass|R.ReadAddressCoef[6]~DUPLICATE_q\ & ((!\TheRxFsk|Lowpass|R.ReadAddressCoef\(2)) # (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(0))))) # (\TheRxFsk|Lowpass|R.ReadAddressCoef\(3) & 
-- (!\TheRxFsk|Lowpass|R.ReadAddressCoef\(2) & ((\TheRxFsk|Lowpass|R.ReadAddressCoef[6]~DUPLICATE_q\)))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1010100001000100101010000100010010001000011000101000100001100010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(3),
	datab => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(2),
	datac => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(0),
	datad => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef[6]~DUPLICATE_q\,
	dataf => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(1),
	combout => \TheRxFsk|Lowpass|CoefMemory~7_combout\);

-- Location: LABCELL_X29_Y67_N12
\TheRxFsk|Lowpass|CoefMemory~8\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|CoefMemory~8_combout\ = ( \TheRxFsk|Lowpass|CoefMemory~7_combout\ & ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(4) & ( !\TheRxFsk|Lowpass|R.ReadAddressCoef\(5) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(5),
	datae => \TheRxFsk|Lowpass|ALT_INV_CoefMemory~7_combout\,
	dataf => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressCoef\(4),
	combout => \TheRxFsk|Lowpass|CoefMemory~8_combout\);

-- Location: M10K_X26_Y65_N0
\TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a0\ : cyclonev_ram_block
-- pragma translate_off
GENERIC MAP (
	mem_init4 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	mem_init3 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	mem_init2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001E00042FFFEDFFFF4FFFE600FFF000160001BFF003FFFE5FFFDE00FF90001E00028FF009FFFDD00FD000FF200026FF038FF013FFFD600FBE00FE70002CFF04BFF02000FD000FAA00FD8FF031FF061FF03100FCD00F9400FC4FF034FF078FF04700FCC00F7CFFFACFF032FF0900006200FCF00F64FFF8FFF02DFF0A70008100FD8FFF4DF",
	mem_init1 => "FF6EFF021000BD000A400FE6FFF38FFF49FF010000D1000CA00FFAFFF27FFF2200FFA000E0000F2FF014FEF1AFFEFA00FDC010EA0011AFF034FEF13FFED201FB9010EDFF140FE05AFFF1400EAD01F91000E9FF164FE084FFF1C01E8B01F66FF0DDFE184FE0B000F2B01E6F00F38FF0C9FE19DFF0DF01F4301E5900F0AFE0AEFE1AE0010D01F6201E4BFFEDDFE08CFF1B80113801F8700E47FEEB3FE065001B80116001FB0FFE4BFEE8EFE039001AF0118200FDDFEE59FEE70FF00B0119C0119CFF00BFEE70FEE5900FDD01182001AFFE039FEE8EFFE4B01FB001160001B8FE065FEEB300E4701F8701138FF1B8FE08CFFEDD01E4B01F620010DFE1AEFE0AE00F",
	mem_init0 => "0A01E5901F43FF0DFFE19DFF0C900F3801E6F00F2BFE0B0FE184FF0DD01F6601E8BFFF1CFE084FF164000E901F9100EADFFF14FE05AFF140010ED01FB9FFED2FEF13FF0340011A010EA00FDCFFEFAFEF1AFF014000F2000E000FFAFFF22FFF2700FFA000CA000D1FF010FFF49FFF3800FE6000A4000BDFF021FFF6EFFF4D00FD800081FF0A7FF02DFFF8F00F6400FCF00062FF090FF032FFFAC00F7C00FCCFF047FF078FF03400FC400F9400FCDFF031FF061FF03100FD800FAA00FD0FF020FF04B0002C00FE700FBEFFFD6FF013FF0380002600FF200FD0FFFDDFF009000280001E00FF9FFFDEFFFE5FF0030001B0001600FFFFFFE6FFFF4FFFED000420001E",
	data_interleave_offset_in_bits => 1,
	data_interleave_width_in_bits => 1,
	init_file => "db/TbdRxFskBasic.ram1_DspFir_da6daf96.hdl.mif",
	init_file_layout => "port_a",
	logical_ram_name => "RxFsk:TheRxFsk|DspFir:\Bandpasses:4:Bandpass0|altsyncram:CoefMemory_rtl_0|altsyncram_gqd1:auto_generated|ALTSYNCRAM",
	operation_mode => "rom",
	port_a_address_clear => "none",
	port_a_address_width => 9,
	port_a_byte_enable_clock => "none",
	port_a_data_out_clear => "none",
	port_a_data_out_clock => "none",
	port_a_data_width => 20,
	port_a_first_address => 0,
	port_a_first_bit_number => 0,
	port_a_last_address => 511,
	port_a_logical_ram_depth => 258,
	port_a_logical_ram_width => 16,
	port_a_read_during_write_mode => "new_data_no_nbe_read",
	port_a_write_enable_clock => "none",
	port_b_address_width => 9,
	port_b_data_width => 20,
	ram_block_type => "M20K")
-- pragma translate_on
PORT MAP (
	portare => VCC,
	clk0 => \iClk~inputCLKENA0_outclk\,
	portaaddr => \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a0_PORTAADDR_bus\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	portadataout => \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a0_PORTADATAOUT_bus\);

-- Location: M10K_X26_Y63_N0
\TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a12\ : cyclonev_ram_block
-- pragma translate_off
GENERIC MAP (
	mem_init4 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	mem_init3 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	mem_init2 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000F0000F0000F0000F0000000000000000000F0000F0000F0000000000000000000F0000F0000F0000000000000000000F0000F0000F0000000000000000000F0000F0000F0000000000000000000F0000F0000F0000000000000000000F0000F0000F0000000000000000000F0000F0000F0000000000000000000F0000F0",
	mem_init1 => "000F0000000000000000000F0000F0000F0000000000000000000F0000F0000F0000F0000000000000000000F0000F0000F0000000000000000000F0000F0000F0000000000000000000F0000F0000F0000000000000000000F0000F0000F0000000000000000000F0000F0000F0000000000000000000F0000F0000F0000000000000000000F0000F0000F0000000000000000000F0000F0000F0000000000000000000F0000F0000F0000000000000000000F0000F0000F000000000000000000000000F0000F0000F0000000000000000000F0000F0000F0000000000000000000F0000F0000F0000000000000000000F0000F0000F000000000000000000",
	mem_init0 => "0F0000F0000F0000000000000000000F0000F0000F0000000000000000000F0000F0000F0000000000000000000F0000F0000F0000000000000000000F0000F0000F0000000000000000000F0000F0000F0000000000000000000F0000F0000F0000F0000000000000000000F0000F0000F0000000000000000000F0000F0000F0000000000000000000F0000F0000F0000000000000000000F0000F0000F0000000000000000000F0000F0000F0000000000000000000F0000F0000F0000000000000000000F0000F0000F0000000000000000000F0000F0000F0000000000000000000F0000F0000F0000000000000000000F0000F0000F0000F0000000000",
	data_interleave_offset_in_bits => 1,
	data_interleave_width_in_bits => 1,
	init_file => "db/TbdRxFskBasic.ram1_DspFir_da6daf96.hdl.mif",
	init_file_layout => "port_a",
	logical_ram_name => "RxFsk:TheRxFsk|DspFir:\Bandpasses:4:Bandpass0|altsyncram:CoefMemory_rtl_0|altsyncram_gqd1:auto_generated|ALTSYNCRAM",
	operation_mode => "rom",
	port_a_address_clear => "none",
	port_a_address_width => 9,
	port_a_byte_enable_clock => "none",
	port_a_data_out_clear => "none",
	port_a_data_out_clock => "none",
	port_a_data_width => 20,
	port_a_first_address => 0,
	port_a_first_bit_number => 12,
	port_a_last_address => 511,
	port_a_logical_ram_depth => 258,
	port_a_logical_ram_width => 16,
	port_a_read_during_write_mode => "new_data_no_nbe_read",
	port_a_write_enable_clock => "none",
	port_b_address_width => 9,
	port_b_data_width => 20,
	ram_block_type => "M20K")
-- pragma translate_on
PORT MAP (
	portare => VCC,
	clk0 => \iClk~inputCLKENA0_outclk\,
	portaaddr => \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a12_PORTAADDR_bus\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	portadataout => \TheRxFsk|Bandpasses:4:Bandpass0|CoefMemory_rtl_0|auto_generated|ram_block1a12_PORTADATAOUT_bus\);

-- Location: IOIBUF_X8_Y81_N1
\iADCdat~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_iADCdat,
	o => \iADCdat~input_o\);

-- Location: LABCELL_X12_Y63_N57
\TheI2sToPar|Decoder0~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheI2sToPar|Decoder0~0_combout\ = ( !\TheI2sToPar|BclkDlyd~q\ & ( (\GenClks|BMclk~q\ & (!\TheI2sToPar|AudioBitCtr\(4) & (!\TheI2sToPar|AudioBitCtr\(3) & \TheI2sToPar|State~q\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001000000000000000100000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \GenClks|ALT_INV_BMclk~q\,
	datab => \TheI2sToPar|ALT_INV_AudioBitCtr\(4),
	datac => \TheI2sToPar|ALT_INV_AudioBitCtr\(3),
	datad => \TheI2sToPar|ALT_INV_State~q\,
	dataf => \TheI2sToPar|ALT_INV_BclkDlyd~q\,
	combout => \TheI2sToPar|Decoder0~0_combout\);

-- Location: LABCELL_X12_Y63_N30
\TheI2sToPar|D[0]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheI2sToPar|D[0]~0_combout\ = ( \TheI2sToPar|Equal0~0_combout\ & ( (!\TheI2sToPar|Decoder0~0_combout\ & ((\TheI2sToPar|D\(0)))) # (\TheI2sToPar|Decoder0~0_combout\ & (\iADCdat~input_o\)) ) ) # ( !\TheI2sToPar|Equal0~0_combout\ & ( \TheI2sToPar|D\(0) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111000011110000111100011101000111010001110100011101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_iADCdat~input_o\,
	datab => \TheI2sToPar|ALT_INV_Decoder0~0_combout\,
	datac => \TheI2sToPar|ALT_INV_D\(0),
	dataf => \TheI2sToPar|ALT_INV_Equal0~0_combout\,
	combout => \TheI2sToPar|D[0]~0_combout\);

-- Location: FF_X15_Y61_N14
\TheI2sToPar|D[0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	asdata => \TheI2sToPar|D[0]~0_combout\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheI2sToPar|D\(0));

-- Location: FF_X15_Y61_N44
\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-15]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	asdata => \TheI2sToPar|D\(0),
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-15]~q\);

-- Location: LABCELL_X13_Y62_N33
\TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[0]~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[0]~1_combout\ = ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(0) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111111111111000000000000000011111111111111110000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.WriteAddress\(0),
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[0]~1_combout\);

-- Location: LABCELL_X13_Y65_N21
\TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[0]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[0]~0_combout\ = ( \TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~q\ & ( (\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~1_combout\ & \TheRxFsk|Bandpasses:11:Bandpass1|Equal1~0_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000001010000010100000000000000000000010100000101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:11:Bandpass1|ALT_INV_Equal1~1_combout\,
	datac => \TheRxFsk|Bandpasses:11:Bandpass1|ALT_INV_Equal1~0_combout\,
	datae => \TheRxFsk|Bandpasses:0:Bandpass0|ALT_INV_R.AddressState~q\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[0]~0_combout\);

-- Location: FF_X13_Y62_N35
\TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[0]~1_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	ena => \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[0]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(0));

-- Location: LABCELL_X13_Y62_N54
\TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[0]~_wirecell\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[0]~_wirecell_combout\ = !\TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(0)

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1010101010101010101010101010101010101010101010101010101010101010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.WriteAddress\(0),
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[0]~_wirecell_combout\);

-- Location: LABCELL_X13_Y62_N0
\TheRxFsk|Bandpasses:4:Bandpass0|Add1~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add1~2\ = CARRY(( !\TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(0) ) + ( VCC ) + ( !VCC ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000000000001111000011110000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.WriteAddress\(0),
	cin => GND,
	cout => \TheRxFsk|Bandpasses:4:Bandpass0|Add1~2\);

-- Location: LABCELL_X13_Y62_N3
\TheRxFsk|Bandpasses:4:Bandpass0|Add1~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add1~5_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(1) ) + ( VCC ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add1~2\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add1~6\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(1) ) + ( VCC ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add1~2\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.WriteAddress\(1),
	cin => \TheRxFsk|Bandpasses:4:Bandpass0|Add1~2\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass0|Add1~5_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass0|Add1~6\);

-- Location: LABCELL_X13_Y62_N6
\TheRxFsk|Bandpasses:4:Bandpass0|Add1~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add1~9_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(2) ) + ( VCC ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add1~6\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add1~10\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(2) ) + ( VCC ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add1~6\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.WriteAddress\(2),
	cin => \TheRxFsk|Bandpasses:4:Bandpass0|Add1~6\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass0|Add1~9_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass0|Add1~10\);

-- Location: FF_X13_Y62_N8
\TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|Add1~9_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:4:Bandpass0|Equal2~1_combout\,
	ena => \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[0]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(2));

-- Location: LABCELL_X13_Y62_N9
\TheRxFsk|Bandpasses:4:Bandpass0|Add1~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add1~13_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(3) ) + ( VCC ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add1~10\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add1~14\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(3) ) + ( VCC ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add1~10\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.WriteAddress\(3),
	cin => \TheRxFsk|Bandpasses:4:Bandpass0|Add1~10\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass0|Add1~13_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass0|Add1~14\);

-- Location: FF_X13_Y62_N10
\TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|Add1~13_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:4:Bandpass0|Equal2~1_combout\,
	ena => \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[0]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(3));

-- Location: LABCELL_X13_Y62_N12
\TheRxFsk|Bandpasses:4:Bandpass0|Add1~17\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add1~17_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(4) ) + ( VCC ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add1~14\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add1~18\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(4) ) + ( VCC ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add1~14\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.WriteAddress\(4),
	cin => \TheRxFsk|Bandpasses:4:Bandpass0|Add1~14\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass0|Add1~17_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass0|Add1~18\);

-- Location: FF_X13_Y62_N13
\TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|Add1~17_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:4:Bandpass0|Equal2~1_combout\,
	ena => \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[0]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(4));

-- Location: LABCELL_X13_Y62_N15
\TheRxFsk|Bandpasses:4:Bandpass0|Add1~21\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add1~21_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(5) ) + ( VCC ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add1~18\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add1~22\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(5) ) + ( VCC ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add1~18\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.WriteAddress\(5),
	cin => \TheRxFsk|Bandpasses:4:Bandpass0|Add1~18\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass0|Add1~21_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass0|Add1~22\);

-- Location: FF_X13_Y62_N16
\TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|Add1~21_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:4:Bandpass0|Equal2~1_combout\,
	ena => \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[0]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(5));

-- Location: LABCELL_X13_Y62_N18
\TheRxFsk|Bandpasses:4:Bandpass0|Add1~25\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add1~25_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(6) ) + ( VCC ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add1~22\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add1~26\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(6) ) + ( VCC ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add1~22\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.WriteAddress\(6),
	cin => \TheRxFsk|Bandpasses:4:Bandpass0|Add1~22\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass0|Add1~25_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass0|Add1~26\);

-- Location: FF_X13_Y62_N19
\TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[6]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|Add1~25_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:4:Bandpass0|Equal2~1_combout\,
	ena => \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[0]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(6));

-- Location: LABCELL_X13_Y62_N21
\TheRxFsk|Bandpasses:4:Bandpass0|Add1~29\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add1~29_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(7) ) + ( VCC ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add1~26\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add1~30\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(7) ) + ( VCC ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add1~26\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.WriteAddress\(7),
	cin => \TheRxFsk|Bandpasses:4:Bandpass0|Add1~26\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass0|Add1~29_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass0|Add1~30\);

-- Location: FF_X13_Y62_N23
\TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[7]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|Add1~29_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:4:Bandpass0|Equal2~1_combout\,
	ena => \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[0]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(7));

-- Location: LABCELL_X13_Y62_N24
\TheRxFsk|Bandpasses:4:Bandpass0|Add1~33\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add1~33_sumout\ = SUM(( !\TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(8) ) + ( VCC ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add1~30\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000000000001100110011001100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.WriteAddress\(8),
	cin => \TheRxFsk|Bandpasses:4:Bandpass0|Add1~30\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass0|Add1~33_sumout\);

-- Location: LABCELL_X13_Y62_N51
\TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[8]~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[8]~2_combout\ = ( !\TheRxFsk|Bandpasses:4:Bandpass0|Add1~33_sumout\ )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111111111111111111111111111100000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add1~33_sumout\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[8]~2_combout\);

-- Location: FF_X13_Y62_N52
\TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[8]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[8]~2_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	ena => \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[0]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(8));

-- Location: LABCELL_X13_Y62_N42
\TheRxFsk|Bandpasses:4:Bandpass0|Equal2~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Equal2~0_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(8) & ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(2) & ( (!\TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(3) & 
-- (!\TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(1) & \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(0))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000010000000100000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.WriteAddress\(3),
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.WriteAddress\(1),
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.WriteAddress\(0),
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.WriteAddress\(8),
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.WriteAddress\(2),
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|Equal2~0_combout\);

-- Location: LABCELL_X13_Y62_N36
\TheRxFsk|Bandpasses:4:Bandpass0|Equal2~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Equal2~1_combout\ = ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(6) & ( (!\TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(5) & (\TheRxFsk|Bandpasses:4:Bandpass0|Equal2~0_combout\ & 
-- (!\TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(7) & !\TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(4)))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0010000000000000001000000000000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.WriteAddress\(5),
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Equal2~0_combout\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.WriteAddress\(7),
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.WriteAddress\(4),
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.WriteAddress\(6),
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|Equal2~1_combout\);

-- Location: FF_X13_Y62_N4
\TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|Add1~5_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:4:Bandpass0|Equal2~1_combout\,
	ena => \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[0]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(1));

-- Location: FF_X13_Y62_N17
\TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[5]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|Add1~21_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:4:Bandpass0|Equal2~1_combout\,
	ena => \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[0]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[5]~DUPLICATE_q\);

-- Location: LABCELL_X13_Y62_N39
\TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[8]~_wirecell\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[8]~_wirecell_combout\ = !\TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress\(8)

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111000011110000111100001111000011110000111100001111000011110000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.WriteAddress\(8),
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|R.WriteAddress[8]~_wirecell_combout\);

-- Location: LABCELL_X13_Y65_N30
\TheRxFsk|Bandpasses:4:Bandpass0|Add0~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add0~1_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(0) ) + ( VCC ) + ( !VCC ))
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add0~2\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(0) ) + ( VCC ) + ( !VCC ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.ReadAddressSample\(0),
	cin => GND,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass0|Add0~1_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass0|Add0~2\);

-- Location: FF_X13_Y65_N31
\TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample[0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|Add0~1_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	ena => \TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(0));

-- Location: LABCELL_X13_Y65_N33
\TheRxFsk|Bandpasses:4:Bandpass0|Add0~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add0~5_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(1) ) + ( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add0~2\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add0~6\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(1) ) + ( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add0~2\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.ReadAddressSample\(1),
	cin => \TheRxFsk|Bandpasses:4:Bandpass0|Add0~2\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass0|Add0~5_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass0|Add0~6\);

-- Location: LABCELL_X13_Y65_N36
\TheRxFsk|Bandpasses:4:Bandpass0|Add0~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add0~9_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(2) ) + ( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add0~6\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add0~10\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(2) ) + ( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add0~6\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.ReadAddressSample\(2),
	cin => \TheRxFsk|Bandpasses:4:Bandpass0|Add0~6\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass0|Add0~9_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass0|Add0~10\);

-- Location: FF_X13_Y65_N37
\TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample[2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|Add0~9_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	ena => \TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(2));

-- Location: LABCELL_X13_Y65_N39
\TheRxFsk|Bandpasses:4:Bandpass0|Add0~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add0~13_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(3) ) + ( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add0~10\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add0~14\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(3) ) + ( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add0~10\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.ReadAddressSample\(3),
	cin => \TheRxFsk|Bandpasses:4:Bandpass0|Add0~10\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass0|Add0~13_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass0|Add0~14\);

-- Location: FF_X13_Y65_N41
\TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample[3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|Add0~13_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	ena => \TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(3));

-- Location: LABCELL_X13_Y65_N42
\TheRxFsk|Bandpasses:4:Bandpass0|Add0~17\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add0~17_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(4) ) + ( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add0~14\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add0~18\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(4) ) + ( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add0~14\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.ReadAddressSample\(4),
	cin => \TheRxFsk|Bandpasses:4:Bandpass0|Add0~14\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass0|Add0~17_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass0|Add0~18\);

-- Location: FF_X13_Y65_N43
\TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample[4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|Add0~17_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	ena => \TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(4));

-- Location: LABCELL_X13_Y65_N45
\TheRxFsk|Bandpasses:4:Bandpass0|Add0~21\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add0~21_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(5) ) + ( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add0~18\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add0~22\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(5) ) + ( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add0~18\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.ReadAddressSample\(5),
	cin => \TheRxFsk|Bandpasses:4:Bandpass0|Add0~18\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass0|Add0~21_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass0|Add0~22\);

-- Location: FF_X13_Y65_N46
\TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample[5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|Add0~21_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	ena => \TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(5));

-- Location: LABCELL_X13_Y65_N48
\TheRxFsk|Bandpasses:4:Bandpass0|Add0~25\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add0~25_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(6) ) + ( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add0~22\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add0~26\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(6) ) + ( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add0~22\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.ReadAddressSample\(6),
	cin => \TheRxFsk|Bandpasses:4:Bandpass0|Add0~22\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass0|Add0~25_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass0|Add0~26\);

-- Location: FF_X13_Y65_N49
\TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample[6]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|Add0~25_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	ena => \TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(6));

-- Location: LABCELL_X13_Y65_N51
\TheRxFsk|Bandpasses:4:Bandpass0|Add0~29\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add0~29_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(7) ) + ( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add0~26\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add0~30\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(7) ) + ( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add0~26\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.ReadAddressSample\(7),
	cin => \TheRxFsk|Bandpasses:4:Bandpass0|Add0~26\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass0|Add0~29_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass0|Add0~30\);

-- Location: FF_X13_Y65_N53
\TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample[7]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|Add0~29_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	ena => \TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(7));

-- Location: LABCELL_X13_Y65_N54
\TheRxFsk|Bandpasses:4:Bandpass0|Add0~33\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add0~33_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(8) ) + ( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add0~30\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.ReadAddressSample\(8),
	cin => \TheRxFsk|Bandpasses:4:Bandpass0|Add0~30\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass0|Add0~33_sumout\);

-- Location: LABCELL_X13_Y65_N27
\TheRxFsk|Bandpasses:4:Bandpass0|NextR~7\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|NextR~7_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(1) & ( \TheRxFsk|Bandpasses:4:Bandpass0|Add0~33_sumout\ ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(1) & ( 
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add0~33_sumout\ & ( (!\TheRxFsk|Bandpasses:4:Bandpass0|Equal0~0_combout\) # (((!\TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(0)) # (\TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(2))) # 
-- (\TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(3))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111101111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Equal0~0_combout\,
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.ReadAddressSample\(3),
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.ReadAddressSample\(2),
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.ReadAddressSample\(0),
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.ReadAddressSample\(1),
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add0~33_sumout\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|NextR~7_combout\);

-- Location: FF_X13_Y65_N28
\TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample[8]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|NextR~7_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	ena => \TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(8));

-- Location: LABCELL_X13_Y65_N0
\TheRxFsk|Bandpasses:4:Bandpass0|Equal0~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Equal0~0_combout\ = ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(5) & ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(7) & ( (!\TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(6) & 
-- (\TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(8) & !\TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(4))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0010000000100000000000000000000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.ReadAddressSample\(6),
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.ReadAddressSample\(8),
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.ReadAddressSample\(4),
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.ReadAddressSample\(5),
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.ReadAddressSample\(7),
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|Equal0~0_combout\);

-- Location: LABCELL_X13_Y65_N24
\TheRxFsk|Bandpasses:4:Bandpass0|NextR~6\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|NextR~6_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(1) & ( \TheRxFsk|Bandpasses:4:Bandpass0|Add0~5_sumout\ ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(1) & ( 
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add0~5_sumout\ & ( (!\TheRxFsk|Bandpasses:4:Bandpass0|Equal0~0_combout\) # (((!\TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(0)) # (\TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(2))) # 
-- (\TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(3))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111011111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Equal0~0_combout\,
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.ReadAddressSample\(3),
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.ReadAddressSample\(0),
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.ReadAddressSample\(2),
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.ReadAddressSample\(1),
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add0~5_sumout\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|NextR~6_combout\);

-- Location: FF_X13_Y65_N25
\TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample[1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|NextR~6_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	ena => \TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|R.ReadAddressSample\(1));

-- Location: LABCELL_X12_Y63_N21
\TheI2sToPar|Decoder0~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheI2sToPar|Decoder0~4_combout\ = ( \TheI2sToPar|AudioBitCtr\(0) & ( !\TheI2sToPar|AudioBitCtr\(3) & ( (\GenClks|BMclk~q\ & (!\TheI2sToPar|AudioBitCtr\(4) & (!\TheI2sToPar|BclkDlyd~q\ & \TheI2sToPar|State~q\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000100000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \GenClks|ALT_INV_BMclk~q\,
	datab => \TheI2sToPar|ALT_INV_AudioBitCtr\(4),
	datac => \TheI2sToPar|ALT_INV_BclkDlyd~q\,
	datad => \TheI2sToPar|ALT_INV_State~q\,
	datae => \TheI2sToPar|ALT_INV_AudioBitCtr\(0),
	dataf => \TheI2sToPar|ALT_INV_AudioBitCtr\(3),
	combout => \TheI2sToPar|Decoder0~4_combout\);

-- Location: MLABCELL_X15_Y63_N0
\TheI2sToPar|D[1]~8\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheI2sToPar|D[1]~8_combout\ = ( \TheI2sToPar|AudioBitCtr[2]~DUPLICATE_q\ & ( \TheI2sToPar|D\(1) ) ) # ( !\TheI2sToPar|AudioBitCtr[2]~DUPLICATE_q\ & ( (!\TheI2sToPar|AudioBitCtr\(1) & ((!\TheI2sToPar|Decoder0~4_combout\ & ((\TheI2sToPar|D\(1)))) # 
-- (\TheI2sToPar|Decoder0~4_combout\ & (\iADCdat~input_o\)))) # (\TheI2sToPar|AudioBitCtr\(1) & (((\TheI2sToPar|D\(1))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010011110111000001001111011100000000111111110000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_iADCdat~input_o\,
	datab => \TheI2sToPar|ALT_INV_AudioBitCtr\(1),
	datac => \TheI2sToPar|ALT_INV_Decoder0~4_combout\,
	datad => \TheI2sToPar|ALT_INV_D\(1),
	dataf => \TheI2sToPar|ALT_INV_AudioBitCtr[2]~DUPLICATE_q\,
	combout => \TheI2sToPar|D[1]~8_combout\);

-- Location: FF_X15_Y63_N8
\TheI2sToPar|D[1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	asdata => \TheI2sToPar|D[1]~8_combout\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheI2sToPar|D\(1));

-- Location: LABCELL_X12_Y63_N36
\TheI2sToPar|D[2]~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheI2sToPar|D[2]~2_combout\ = ( \TheI2sToPar|AudioBitCtr[1]~DUPLICATE_q\ & ( \TheI2sToPar|AudioBitCtr\(2) & ( \TheI2sToPar|D\(2) ) ) ) # ( !\TheI2sToPar|AudioBitCtr[1]~DUPLICATE_q\ & ( \TheI2sToPar|AudioBitCtr\(2) & ( \TheI2sToPar|D\(2) ) ) ) # ( 
-- \TheI2sToPar|AudioBitCtr[1]~DUPLICATE_q\ & ( !\TheI2sToPar|AudioBitCtr\(2) & ( (!\TheI2sToPar|Decoder0~0_combout\ & (\TheI2sToPar|D\(2))) # (\TheI2sToPar|Decoder0~0_combout\ & ((!\TheI2sToPar|AudioBitCtr\(0) & ((\iADCdat~input_o\))) # 
-- (\TheI2sToPar|AudioBitCtr\(0) & (\TheI2sToPar|D\(2))))) ) ) ) # ( !\TheI2sToPar|AudioBitCtr[1]~DUPLICATE_q\ & ( !\TheI2sToPar|AudioBitCtr\(2) & ( \TheI2sToPar|D\(2) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010101010101010001110101010101010101010101010101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheI2sToPar|ALT_INV_D\(2),
	datab => \TheI2sToPar|ALT_INV_Decoder0~0_combout\,
	datac => \ALT_INV_iADCdat~input_o\,
	datad => \TheI2sToPar|ALT_INV_AudioBitCtr\(0),
	datae => \TheI2sToPar|ALT_INV_AudioBitCtr[1]~DUPLICATE_q\,
	dataf => \TheI2sToPar|ALT_INV_AudioBitCtr\(2),
	combout => \TheI2sToPar|D[2]~2_combout\);

-- Location: FF_X13_Y63_N11
\TheI2sToPar|D[2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	asdata => \TheI2sToPar|D[2]~2_combout\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheI2sToPar|D\(2));

-- Location: LABCELL_X16_Y63_N36
\TheI2sToPar|D[3]~10\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheI2sToPar|D[3]~10_combout\ = ( \TheI2sToPar|AudioBitCtr[2]~DUPLICATE_q\ & ( \TheI2sToPar|D\(3) ) ) # ( !\TheI2sToPar|AudioBitCtr[2]~DUPLICATE_q\ & ( (!\TheI2sToPar|Decoder0~4_combout\ & (((\TheI2sToPar|D\(3))))) # (\TheI2sToPar|Decoder0~4_combout\ & 
-- ((!\TheI2sToPar|AudioBitCtr[1]~DUPLICATE_q\ & ((\TheI2sToPar|D\(3)))) # (\TheI2sToPar|AudioBitCtr[1]~DUPLICATE_q\ & (\iADCdat~input_o\)))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001100110101001100110011010100110011001100110011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_iADCdat~input_o\,
	datab => \TheI2sToPar|ALT_INV_D\(3),
	datac => \TheI2sToPar|ALT_INV_Decoder0~4_combout\,
	datad => \TheI2sToPar|ALT_INV_AudioBitCtr[1]~DUPLICATE_q\,
	dataf => \TheI2sToPar|ALT_INV_AudioBitCtr[2]~DUPLICATE_q\,
	combout => \TheI2sToPar|D[3]~10_combout\);

-- Location: FF_X15_Y63_N38
\TheI2sToPar|D[3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	asdata => \TheI2sToPar|D[3]~10_combout\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheI2sToPar|D\(3));

-- Location: MLABCELL_X15_Y63_N3
\TheI2sToPar|Equal0~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheI2sToPar|Equal0~2_combout\ = (!\TheI2sToPar|AudioBitCtr\(1) & !\TheI2sToPar|AudioBitCtr\(0))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1100000011000000110000001100000011000000110000001100000011000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheI2sToPar|ALT_INV_AudioBitCtr\(1),
	datac => \TheI2sToPar|ALT_INV_AudioBitCtr\(0),
	combout => \TheI2sToPar|Equal0~2_combout\);

-- Location: MLABCELL_X15_Y63_N45
\TheI2sToPar|D[4]~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheI2sToPar|D[4]~4_combout\ = ( \TheI2sToPar|Equal0~2_combout\ & ( \TheI2sToPar|AudioBitCtr[2]~DUPLICATE_q\ & ( (!\TheI2sToPar|Decoder0~0_combout\ & (\TheI2sToPar|D\(4))) # (\TheI2sToPar|Decoder0~0_combout\ & ((\iADCdat~input_o\))) ) ) ) # ( 
-- !\TheI2sToPar|Equal0~2_combout\ & ( \TheI2sToPar|AudioBitCtr[2]~DUPLICATE_q\ & ( \TheI2sToPar|D\(4) ) ) ) # ( \TheI2sToPar|Equal0~2_combout\ & ( !\TheI2sToPar|AudioBitCtr[2]~DUPLICATE_q\ & ( \TheI2sToPar|D\(4) ) ) ) # ( !\TheI2sToPar|Equal0~2_combout\ & ( 
-- !\TheI2sToPar|AudioBitCtr[2]~DUPLICATE_q\ & ( \TheI2sToPar|D\(4) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010101010101010101010101010101010101010101010101001101010011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheI2sToPar|ALT_INV_D\(4),
	datab => \ALT_INV_iADCdat~input_o\,
	datac => \TheI2sToPar|ALT_INV_Decoder0~0_combout\,
	datae => \TheI2sToPar|ALT_INV_Equal0~2_combout\,
	dataf => \TheI2sToPar|ALT_INV_AudioBitCtr[2]~DUPLICATE_q\,
	combout => \TheI2sToPar|D[4]~4_combout\);

-- Location: FF_X15_Y63_N50
\TheI2sToPar|D[4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	asdata => \TheI2sToPar|D[4]~4_combout\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheI2sToPar|D\(4));

-- Location: MLABCELL_X15_Y63_N48
\TheI2sToPar|D[5]~12\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheI2sToPar|D[5]~12_combout\ = ( \TheI2sToPar|AudioBitCtr[2]~DUPLICATE_q\ & ( (!\TheI2sToPar|AudioBitCtr\(1) & ((!\TheI2sToPar|Decoder0~4_combout\ & (\TheI2sToPar|D\(5))) # (\TheI2sToPar|Decoder0~4_combout\ & ((\iADCdat~input_o\))))) # 
-- (\TheI2sToPar|AudioBitCtr\(1) & (\TheI2sToPar|D\(5))) ) ) # ( !\TheI2sToPar|AudioBitCtr[2]~DUPLICATE_q\ & ( \TheI2sToPar|D\(5) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010101010101010101010101010101010001010111010101000101011101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheI2sToPar|ALT_INV_D\(5),
	datab => \TheI2sToPar|ALT_INV_AudioBitCtr\(1),
	datac => \TheI2sToPar|ALT_INV_Decoder0~4_combout\,
	datad => \ALT_INV_iADCdat~input_o\,
	dataf => \TheI2sToPar|ALT_INV_AudioBitCtr[2]~DUPLICATE_q\,
	combout => \TheI2sToPar|D[5]~12_combout\);

-- Location: FF_X13_Y62_N59
\TheI2sToPar|D[5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	asdata => \TheI2sToPar|D[5]~12_combout\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheI2sToPar|D\(5));

-- Location: LABCELL_X12_Y63_N3
\TheI2sToPar|Decoder0~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheI2sToPar|Decoder0~3_combout\ = ( \TheI2sToPar|AudioBitCtr\(2) & ( \TheI2sToPar|AudioBitCtr[1]~DUPLICATE_q\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000111111110000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \TheI2sToPar|ALT_INV_AudioBitCtr[1]~DUPLICATE_q\,
	dataf => \TheI2sToPar|ALT_INV_AudioBitCtr\(2),
	combout => \TheI2sToPar|Decoder0~3_combout\);

-- Location: LABCELL_X12_Y63_N33
\TheI2sToPar|D[6]~6\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheI2sToPar|D[6]~6_combout\ = ( \TheI2sToPar|D\(6) & ( ((!\TheI2sToPar|Decoder0~0_combout\) # ((!\TheI2sToPar|Decoder0~3_combout\) # (\TheI2sToPar|AudioBitCtr\(0)))) # (\iADCdat~input_o\) ) ) # ( !\TheI2sToPar|D\(6) & ( (\iADCdat~input_o\ & 
-- (\TheI2sToPar|Decoder0~0_combout\ & (!\TheI2sToPar|AudioBitCtr\(0) & \TheI2sToPar|Decoder0~3_combout\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000010000000000000001000011111111110111111111111111011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_iADCdat~input_o\,
	datab => \TheI2sToPar|ALT_INV_Decoder0~0_combout\,
	datac => \TheI2sToPar|ALT_INV_AudioBitCtr\(0),
	datad => \TheI2sToPar|ALT_INV_Decoder0~3_combout\,
	dataf => \TheI2sToPar|ALT_INV_D\(6),
	combout => \TheI2sToPar|D[6]~6_combout\);

-- Location: FF_X15_Y63_N2
\TheI2sToPar|D[6]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	asdata => \TheI2sToPar|D[6]~6_combout\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheI2sToPar|D\(6));

-- Location: LABCELL_X13_Y64_N12
\TheI2sToPar|D[7]~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheI2sToPar|D[7]~14_combout\ = ( \iADCdat~input_o\ & ( \TheI2sToPar|D\(7) ) ) # ( !\iADCdat~input_o\ & ( \TheI2sToPar|D\(7) & ( (!\TheI2sToPar|Decoder0~3_combout\) # (!\TheI2sToPar|Decoder0~4_combout\) ) ) ) # ( \iADCdat~input_o\ & ( !\TheI2sToPar|D\(7) 
-- & ( (\TheI2sToPar|Decoder0~3_combout\ & \TheI2sToPar|Decoder0~4_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000100010001000111101110111011101111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheI2sToPar|ALT_INV_Decoder0~3_combout\,
	datab => \TheI2sToPar|ALT_INV_Decoder0~4_combout\,
	datae => \ALT_INV_iADCdat~input_o\,
	dataf => \TheI2sToPar|ALT_INV_D\(7),
	combout => \TheI2sToPar|D[7]~14_combout\);

-- Location: FF_X13_Y64_N26
\TheI2sToPar|D[7]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	asdata => \TheI2sToPar|D[7]~14_combout\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheI2sToPar|D\(7));

-- Location: LABCELL_X12_Y63_N18
\TheI2sToPar|Decoder0~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheI2sToPar|Decoder0~1_combout\ = ( \TheI2sToPar|AudioBitCtr\(3) & ( !\TheI2sToPar|AudioBitCtr\(2) & ( (\GenClks|BMclk~q\ & (!\TheI2sToPar|AudioBitCtr\(4) & (\TheI2sToPar|State~q\ & !\TheI2sToPar|BclkDlyd~q\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000001000000000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \GenClks|ALT_INV_BMclk~q\,
	datab => \TheI2sToPar|ALT_INV_AudioBitCtr\(4),
	datac => \TheI2sToPar|ALT_INV_State~q\,
	datad => \TheI2sToPar|ALT_INV_BclkDlyd~q\,
	datae => \TheI2sToPar|ALT_INV_AudioBitCtr\(3),
	dataf => \TheI2sToPar|ALT_INV_AudioBitCtr\(2),
	combout => \TheI2sToPar|Decoder0~1_combout\);

-- Location: MLABCELL_X15_Y63_N24
\TheI2sToPar|D[8]~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheI2sToPar|D[8]~1_combout\ = ( \TheI2sToPar|D\(8) & ( (!\TheI2sToPar|Decoder0~1_combout\) # ((!\TheI2sToPar|Equal0~2_combout\) # (\iADCdat~input_o\)) ) ) # ( !\TheI2sToPar|D\(8) & ( (\TheI2sToPar|Decoder0~1_combout\ & (\iADCdat~input_o\ & 
-- \TheI2sToPar|Equal0~2_combout\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000100000001000000010000000111111011111110111111101111111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheI2sToPar|ALT_INV_Decoder0~1_combout\,
	datab => \ALT_INV_iADCdat~input_o\,
	datac => \TheI2sToPar|ALT_INV_Equal0~2_combout\,
	dataf => \TheI2sToPar|ALT_INV_D\(8),
	combout => \TheI2sToPar|D[8]~1_combout\);

-- Location: FF_X13_Y63_N26
\TheI2sToPar|D[8]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	asdata => \TheI2sToPar|D[8]~1_combout\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheI2sToPar|D\(8));

-- Location: MLABCELL_X15_Y63_N27
\TheI2sToPar|D[9]~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheI2sToPar|D[9]~9_combout\ = ( \TheI2sToPar|AudioBitCtr\(0) & ( (!\TheI2sToPar|Decoder0~1_combout\ & (((\TheI2sToPar|D\(9))))) # (\TheI2sToPar|Decoder0~1_combout\ & ((!\TheI2sToPar|AudioBitCtr\(1) & (\iADCdat~input_o\)) # (\TheI2sToPar|AudioBitCtr\(1) & 
-- ((\TheI2sToPar|D\(9)))))) ) ) # ( !\TheI2sToPar|AudioBitCtr\(0) & ( \TheI2sToPar|D\(9) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011111111000000001111111100010000101111110001000010111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheI2sToPar|ALT_INV_Decoder0~1_combout\,
	datab => \ALT_INV_iADCdat~input_o\,
	datac => \TheI2sToPar|ALT_INV_AudioBitCtr\(1),
	datad => \TheI2sToPar|ALT_INV_D\(9),
	dataf => \TheI2sToPar|ALT_INV_AudioBitCtr\(0),
	combout => \TheI2sToPar|D[9]~9_combout\);

-- Location: FF_X15_Y63_N26
\TheI2sToPar|D[9]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	asdata => \TheI2sToPar|D[9]~9_combout\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheI2sToPar|D\(9));

-- Location: LABCELL_X16_Y63_N24
\TheI2sToPar|D[10]~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheI2sToPar|D[10]~3_combout\ = ( \TheI2sToPar|D\(10) & ( ((!\TheI2sToPar|AudioBitCtr[1]~DUPLICATE_q\) # ((!\TheI2sToPar|Decoder0~1_combout\) # (\iADCdat~input_o\))) # (\TheI2sToPar|AudioBitCtr\(0)) ) ) # ( !\TheI2sToPar|D\(10) & ( 
-- (!\TheI2sToPar|AudioBitCtr\(0) & (\TheI2sToPar|AudioBitCtr[1]~DUPLICATE_q\ & (\iADCdat~input_o\ & \TheI2sToPar|Decoder0~1_combout\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000010000000000000001011111111110111111111111111011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheI2sToPar|ALT_INV_AudioBitCtr\(0),
	datab => \TheI2sToPar|ALT_INV_AudioBitCtr[1]~DUPLICATE_q\,
	datac => \ALT_INV_iADCdat~input_o\,
	datad => \TheI2sToPar|ALT_INV_Decoder0~1_combout\,
	dataf => \TheI2sToPar|ALT_INV_D\(10),
	combout => \TheI2sToPar|D[10]~3_combout\);

-- Location: FF_X15_Y63_N44
\TheI2sToPar|D[10]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	asdata => \TheI2sToPar|D[10]~3_combout\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheI2sToPar|D\(10));

-- Location: LABCELL_X16_Y63_N27
\TheI2sToPar|D[11]~11\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheI2sToPar|D[11]~11_combout\ = ( \iADCdat~input_o\ & ( ((\TheI2sToPar|AudioBitCtr\(0) & (\TheI2sToPar|AudioBitCtr[1]~DUPLICATE_q\ & \TheI2sToPar|Decoder0~1_combout\))) # (\TheI2sToPar|D\(11)) ) ) # ( !\iADCdat~input_o\ & ( (\TheI2sToPar|D\(11) & 
-- ((!\TheI2sToPar|AudioBitCtr\(0)) # ((!\TheI2sToPar|AudioBitCtr[1]~DUPLICATE_q\) # (!\TheI2sToPar|Decoder0~1_combout\)))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001110000011110000111000001111000111110000111100011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheI2sToPar|ALT_INV_AudioBitCtr\(0),
	datab => \TheI2sToPar|ALT_INV_AudioBitCtr[1]~DUPLICATE_q\,
	datac => \TheI2sToPar|ALT_INV_D\(11),
	datad => \TheI2sToPar|ALT_INV_Decoder0~1_combout\,
	dataf => \ALT_INV_iADCdat~input_o\,
	combout => \TheI2sToPar|D[11]~11_combout\);

-- Location: FF_X15_Y63_N59
\TheI2sToPar|D[11]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	asdata => \TheI2sToPar|D[11]~11_combout\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheI2sToPar|D\(11));

-- Location: LABCELL_X12_Y63_N54
\TheI2sToPar|Decoder0~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheI2sToPar|Decoder0~2_combout\ = ( !\TheI2sToPar|BclkDlyd~q\ & ( (\GenClks|BMclk~q\ & (!\TheI2sToPar|AudioBitCtr\(4) & (\TheI2sToPar|State~q\ & \TheI2sToPar|AudioBitCtr\(3)))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000100000000000000010000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \GenClks|ALT_INV_BMclk~q\,
	datab => \TheI2sToPar|ALT_INV_AudioBitCtr\(4),
	datac => \TheI2sToPar|ALT_INV_State~q\,
	datad => \TheI2sToPar|ALT_INV_AudioBitCtr\(3),
	dataf => \TheI2sToPar|ALT_INV_BclkDlyd~q\,
	combout => \TheI2sToPar|Decoder0~2_combout\);

-- Location: LABCELL_X16_Y63_N45
\TheI2sToPar|D[12]~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheI2sToPar|D[12]~5_combout\ = ( \TheI2sToPar|Decoder0~2_combout\ & ( \TheI2sToPar|Equal0~2_combout\ & ( (!\TheI2sToPar|AudioBitCtr[2]~DUPLICATE_q\ & ((\TheI2sToPar|D\(12)))) # (\TheI2sToPar|AudioBitCtr[2]~DUPLICATE_q\ & (\iADCdat~input_o\)) ) ) ) # ( 
-- !\TheI2sToPar|Decoder0~2_combout\ & ( \TheI2sToPar|Equal0~2_combout\ & ( \TheI2sToPar|D\(12) ) ) ) # ( \TheI2sToPar|Decoder0~2_combout\ & ( !\TheI2sToPar|Equal0~2_combout\ & ( \TheI2sToPar|D\(12) ) ) ) # ( !\TheI2sToPar|Decoder0~2_combout\ & ( 
-- !\TheI2sToPar|Equal0~2_combout\ & ( \TheI2sToPar|D\(12) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011111111000000001111111100000000111111110000010111110101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \ALT_INV_iADCdat~input_o\,
	datac => \TheI2sToPar|ALT_INV_AudioBitCtr[2]~DUPLICATE_q\,
	datad => \TheI2sToPar|ALT_INV_D\(12),
	datae => \TheI2sToPar|ALT_INV_Decoder0~2_combout\,
	dataf => \TheI2sToPar|ALT_INV_Equal0~2_combout\,
	combout => \TheI2sToPar|D[12]~5_combout\);

-- Location: FF_X15_Y63_N53
\TheI2sToPar|D[12]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	asdata => \TheI2sToPar|D[12]~5_combout\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheI2sToPar|D\(12));

-- Location: LABCELL_X16_Y63_N54
\TheI2sToPar|D[13]~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheI2sToPar|D[13]~13_combout\ = ( \TheI2sToPar|AudioBitCtr[1]~DUPLICATE_q\ & ( \iADCdat~input_o\ & ( \TheI2sToPar|D\(13) ) ) ) # ( !\TheI2sToPar|AudioBitCtr[1]~DUPLICATE_q\ & ( \iADCdat~input_o\ & ( ((\TheI2sToPar|Decoder0~2_combout\ & 
-- (\TheI2sToPar|AudioBitCtr\(0) & \TheI2sToPar|AudioBitCtr[2]~DUPLICATE_q\))) # (\TheI2sToPar|D\(13)) ) ) ) # ( \TheI2sToPar|AudioBitCtr[1]~DUPLICATE_q\ & ( !\iADCdat~input_o\ & ( \TheI2sToPar|D\(13) ) ) ) # ( !\TheI2sToPar|AudioBitCtr[1]~DUPLICATE_q\ & ( 
-- !\iADCdat~input_o\ & ( (\TheI2sToPar|D\(13) & ((!\TheI2sToPar|Decoder0~2_combout\) # ((!\TheI2sToPar|AudioBitCtr\(0)) # (!\TheI2sToPar|AudioBitCtr[2]~DUPLICATE_q\)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010101010100010101010101010101010101010101110101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheI2sToPar|ALT_INV_D\(13),
	datab => \TheI2sToPar|ALT_INV_Decoder0~2_combout\,
	datac => \TheI2sToPar|ALT_INV_AudioBitCtr\(0),
	datad => \TheI2sToPar|ALT_INV_AudioBitCtr[2]~DUPLICATE_q\,
	datae => \TheI2sToPar|ALT_INV_AudioBitCtr[1]~DUPLICATE_q\,
	dataf => \ALT_INV_iADCdat~input_o\,
	combout => \TheI2sToPar|D[13]~13_combout\);

-- Location: FF_X15_Y63_N41
\TheI2sToPar|D[13]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	asdata => \TheI2sToPar|D[13]~13_combout\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheI2sToPar|D\(13));

-- Location: LABCELL_X12_Y63_N6
\TheI2sToPar|D[14]~7\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheI2sToPar|D[14]~7_combout\ = ( \iADCdat~input_o\ & ( ((\TheI2sToPar|Decoder0~3_combout\ & (!\TheI2sToPar|AudioBitCtr\(0) & \TheI2sToPar|Decoder0~2_combout\))) # (\TheI2sToPar|D\(14)) ) ) # ( !\iADCdat~input_o\ & ( (\TheI2sToPar|D\(14) & 
-- ((!\TheI2sToPar|Decoder0~3_combout\) # ((!\TheI2sToPar|Decoder0~2_combout\) # (\TheI2sToPar|AudioBitCtr\(0))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011111011000000001111101100000100111111110000010011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheI2sToPar|ALT_INV_Decoder0~3_combout\,
	datab => \TheI2sToPar|ALT_INV_AudioBitCtr\(0),
	datac => \TheI2sToPar|ALT_INV_Decoder0~2_combout\,
	datad => \TheI2sToPar|ALT_INV_D\(14),
	dataf => \ALT_INV_iADCdat~input_o\,
	combout => \TheI2sToPar|D[14]~7_combout\);

-- Location: MLABCELL_X15_Y63_N9
\TheI2sToPar|D[14]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheI2sToPar|D[14]~feeder_combout\ = ( \TheI2sToPar|D[14]~7_combout\ )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \TheI2sToPar|ALT_INV_D[14]~7_combout\,
	combout => \TheI2sToPar|D[14]~feeder_combout\);

-- Location: FF_X15_Y63_N11
\TheI2sToPar|D[14]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \TheI2sToPar|D[14]~feeder_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheI2sToPar|D\(14));

-- Location: LABCELL_X12_Y63_N9
\TheI2sToPar|D[15]~15\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheI2sToPar|D[15]~15_combout\ = ( \TheI2sToPar|Decoder0~2_combout\ & ( (!\TheI2sToPar|Decoder0~3_combout\ & (((\TheI2sToPar|D\(15))))) # (\TheI2sToPar|Decoder0~3_combout\ & ((!\TheI2sToPar|AudioBitCtr\(0) & (\TheI2sToPar|D\(15))) # 
-- (\TheI2sToPar|AudioBitCtr\(0) & ((\iADCdat~input_o\))))) ) ) # ( !\TheI2sToPar|Decoder0~2_combout\ & ( \TheI2sToPar|D\(15) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111000011110000111100001110000111110000111000011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheI2sToPar|ALT_INV_Decoder0~3_combout\,
	datab => \TheI2sToPar|ALT_INV_AudioBitCtr\(0),
	datac => \TheI2sToPar|ALT_INV_D\(15),
	datad => \ALT_INV_iADCdat~input_o\,
	dataf => \TheI2sToPar|ALT_INV_Decoder0~2_combout\,
	combout => \TheI2sToPar|D[15]~15_combout\);

-- Location: FF_X13_Y63_N8
\TheI2sToPar|D[15]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	asdata => \TheI2sToPar|D[15]~15_combout\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheI2sToPar|D\(15));

-- Location: M10K_X14_Y64_N0
\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a0\ : cyclonev_ram_block
-- pragma translate_off
GENERIC MAP (
	mem_init4 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	mem_init3 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	mem_init2 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	mem_init1 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	mem_init0 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	data_interleave_offset_in_bits => 1,
	data_interleave_width_in_bits => 1,
	init_file => "db/TbdRxFskBasic.ram0_DspFir_da6daf96.hdl.mif",
	init_file_layout => "port_a",
	logical_ram_name => "RxFsk:TheRxFsk|DspFir:\Bandpasses:4:Bandpass0|altsyncram:SampleMemory_rtl_0|altsyncram_qes1:auto_generated|ALTSYNCRAM",
	mixed_port_feed_through_mode => "old",
	operation_mode => "dual_port",
	port_a_address_clear => "none",
	port_a_address_width => 9,
	port_a_byte_enable_clock => "none",
	port_a_data_out_clear => "none",
	port_a_data_out_clock => "none",
	port_a_data_width => 20,
	port_a_first_address => 0,
	port_a_first_bit_number => 0,
	port_a_last_address => 511,
	port_a_logical_ram_depth => 258,
	port_a_logical_ram_width => 16,
	port_a_read_during_write_mode => "new_data_no_nbe_read",
	port_b_address_clear => "none",
	port_b_address_clock => "clock0",
	port_b_address_width => 9,
	port_b_data_out_clear => "none",
	port_b_data_out_clock => "none",
	port_b_data_width => 20,
	port_b_first_address => 0,
	port_b_first_bit_number => 0,
	port_b_last_address => 511,
	port_b_logical_ram_depth => 258,
	port_b_logical_ram_width => 16,
	port_b_read_during_write_mode => "new_data_no_nbe_read",
	port_b_read_enable_clock => "clock0",
	ram_block_type => "M20K")
-- pragma translate_on
PORT MAP (
	portawe => \TheI2sToPar|ValL~q\,
	portbre => VCC,
	clk0 => \iClk~inputCLKENA0_outclk\,
	portadatain => \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTADATAIN_bus\,
	portaaddr => \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTAADDR_bus\,
	portbaddr => \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBADDR_bus\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	portbdataout => \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\);

-- Location: FF_X17_Y65_N55
\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	asdata => \TheRxFsk|Bandpasses:0:Bandpass0|R.AddressState~q\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\);

-- Location: LABCELL_X16_Y65_N33
\TheRxFsk|Bandpasses:4:Bandpass0|Sample[-15]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-15]~0_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a0~portbdataout\ ) ) # ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-15]~q\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111000011110000111100000000111111110000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-15]~q\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a0~portbdataout\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-15]~0_combout\);

-- Location: FF_X15_Y63_N23
\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-14]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	asdata => \TheI2sToPar|D\(1),
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-14]~q\);

-- Location: LABCELL_X16_Y62_N6
\TheRxFsk|Bandpasses:4:Bandpass0|Sample[-14]~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-14]~1_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a1\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\) # (\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-14]~q\) ) 
-- ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a1\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-14]~q\ & !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001100000000001100110000000000110011111111110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-14]~q\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a1\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-14]~1_combout\);

-- Location: FF_X13_Y63_N20
\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-13]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	asdata => \TheI2sToPar|D\(2),
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-13]~q\);

-- Location: LABCELL_X19_Y63_N33
\TheRxFsk|Bandpasses:4:Bandpass0|Sample[-13]~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-13]~2_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a2\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-13]~q\) # (\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\) ) 
-- ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a2\ & ( (!\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-13]~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000101000001010000010100000101001011111010111110101111101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-13]~q\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a2\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-13]~2_combout\);

-- Location: FF_X15_Y63_N17
\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-12]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	asdata => \TheI2sToPar|D\(3),
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-12]~q\);

-- Location: LABCELL_X18_Y65_N30
\TheRxFsk|Bandpasses:4:Bandpass0|Sample[-12]~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-12]~3_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-12]~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a3\ ) ) # ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-12]~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a3\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ ) ) ) # ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-12]~q\ 
-- & ( !\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a3\ & ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000001111000011111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-12]~q\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a3\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-12]~3_combout\);

-- Location: LABCELL_X16_Y63_N48
\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-11]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-11]~feeder_combout\ = ( \TheI2sToPar|D\(4) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \TheI2sToPar|ALT_INV_D\(4),
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-11]~feeder_combout\);

-- Location: FF_X16_Y63_N49
\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-11]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-11]~feeder_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-11]~q\);

-- Location: LABCELL_X17_Y63_N33
\TheRxFsk|Bandpasses:4:Bandpass0|Sample[-11]~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-11]~4_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-11]~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a4\ ) ) # ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-11]~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a4\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ ) ) ) # ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-11]~q\ 
-- & ( !\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a4\ & ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000101010101010101001010101010101011111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-11]~q\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a4\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-11]~4_combout\);

-- Location: FF_X13_Y62_N28
\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-10]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	asdata => \TheI2sToPar|D\(5),
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-10]~q\);

-- Location: LABCELL_X17_Y63_N36
\TheRxFsk|Bandpasses:4:Bandpass0|Sample[-10]~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-10]~5_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a5\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-10]~q\ ) ) # ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a5\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-10]~q\ & ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ ) ) ) # ( 
-- \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a5\ & ( !\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-10]~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000010101010101010110101010101010101111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a5\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-10]~q\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-10]~5_combout\);

-- Location: FF_X15_Y63_N20
\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-9]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	asdata => \TheI2sToPar|D\(6),
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-9]~q\);

-- Location: LABCELL_X17_Y63_N9
\TheRxFsk|Bandpasses:4:Bandpass0|Sample[-9]~6\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-9]~6_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a6\ ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & 
-- ( \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a6\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-9]~q\ ) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a6\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-9]~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111000000000000000000001111000011111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-9]~q\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a6\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-9]~6_combout\);

-- Location: FF_X13_Y64_N38
\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-8]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	asdata => \TheI2sToPar|D\(7),
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-8]~q\);

-- Location: LABCELL_X13_Y64_N36
\TheRxFsk|Bandpasses:4:Bandpass0|Sample[-8]~7\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-8]~7_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a7\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-8]~q\) # (\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\) ) ) 
-- # ( !\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a7\ & ( (!\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-8]~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011001100000000001100110000110011111111110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-8]~q\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a7\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-8]~7_combout\);

-- Location: FF_X15_Y63_N31
\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-7]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	asdata => \TheI2sToPar|D\(8),
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-7]~q\);

-- Location: LABCELL_X18_Y65_N0
\TheRxFsk|Bandpasses:4:Bandpass0|Sample[-7]~8\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-7]~8_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a8\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\) # (\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-7]~q\) ) ) 
-- # ( !\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a8\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-7]~q\ & !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101000001010000010111110101111101010000010100000101111101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-7]~q\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a8\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-7]~8_combout\);

-- Location: FF_X15_Y63_N35
\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-6]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	asdata => \TheI2sToPar|D\(9),
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-6]~q\);

-- Location: MLABCELL_X15_Y65_N24
\TheRxFsk|Bandpasses:4:Bandpass0|Sample[-6]~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-6]~9_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a9\ ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & 
-- ( \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a9\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-6]~q\ ) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a9\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-6]~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001100110011000000000000000000110011001100111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-6]~q\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a9\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-6]~9_combout\);

-- Location: LABCELL_X16_Y63_N51
\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-5]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-5]~feeder_combout\ = ( \TheI2sToPar|D\(10) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \TheI2sToPar|ALT_INV_D\(10),
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-5]~feeder_combout\);

-- Location: FF_X16_Y63_N52
\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-5]~feeder_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-5]~q\);

-- Location: LABCELL_X18_Y65_N54
\TheRxFsk|Bandpasses:4:Bandpass0|Sample[-5]~10\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-5]~10_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a10\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-5]~q\ ) ) # ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a10\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-5]~q\ & ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ ) ) ) # ( 
-- \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a10\ & ( !\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-5]~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000011110000111111110000111100001111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a10\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-5]~q\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-5]~10_combout\);

-- Location: LABCELL_X16_Y63_N0
\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-4]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-4]~feeder_combout\ = ( \TheI2sToPar|D\(11) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \TheI2sToPar|ALT_INV_D\(11),
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-4]~feeder_combout\);

-- Location: FF_X16_Y63_N1
\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-4]~feeder_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-4]~q\);

-- Location: MLABCELL_X15_Y65_N54
\TheRxFsk|Bandpasses:4:Bandpass0|Sample[-4]~11\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-4]~11_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a11\ ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ 
-- & ( \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a11\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-4]~q\ ) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a11\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-4]~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111000000000000000000001111000011111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-4]~q\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a11\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-4]~11_combout\);

-- Location: FF_X15_Y63_N14
\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	asdata => \TheI2sToPar|D\(12),
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-3]~q\);

-- Location: M10K_X14_Y65_N0
\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a12\ : cyclonev_ram_block
-- pragma translate_off
GENERIC MAP (
	mem_init4 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	mem_init3 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	mem_init2 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	mem_init1 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	mem_init0 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	data_interleave_offset_in_bits => 1,
	data_interleave_width_in_bits => 1,
	init_file => "db/TbdRxFskBasic.ram0_DspFir_da6daf96.hdl.mif",
	init_file_layout => "port_a",
	logical_ram_name => "RxFsk:TheRxFsk|DspFir:\Bandpasses:4:Bandpass0|altsyncram:SampleMemory_rtl_0|altsyncram_qes1:auto_generated|ALTSYNCRAM",
	mixed_port_feed_through_mode => "old",
	operation_mode => "dual_port",
	port_a_address_clear => "none",
	port_a_address_width => 9,
	port_a_byte_enable_clock => "none",
	port_a_data_out_clear => "none",
	port_a_data_out_clock => "none",
	port_a_data_width => 20,
	port_a_first_address => 0,
	port_a_first_bit_number => 12,
	port_a_last_address => 511,
	port_a_logical_ram_depth => 258,
	port_a_logical_ram_width => 16,
	port_a_read_during_write_mode => "new_data_no_nbe_read",
	port_b_address_clear => "none",
	port_b_address_clock => "clock0",
	port_b_address_width => 9,
	port_b_data_out_clear => "none",
	port_b_data_out_clock => "none",
	port_b_data_width => 20,
	port_b_first_address => 0,
	port_b_first_bit_number => 12,
	port_b_last_address => 511,
	port_b_logical_ram_depth => 258,
	port_b_logical_ram_width => 16,
	port_b_read_during_write_mode => "new_data_no_nbe_read",
	port_b_read_enable_clock => "clock0",
	ram_block_type => "M20K")
-- pragma translate_on
PORT MAP (
	portawe => \TheI2sToPar|ValL~q\,
	portbre => VCC,
	clk0 => \iClk~inputCLKENA0_outclk\,
	portadatain => \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a12_PORTADATAIN_bus\,
	portaaddr => \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a12_PORTAADDR_bus\,
	portbaddr => \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a12_PORTBADDR_bus\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	portbdataout => \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a12_PORTBDATAOUT_bus\);

-- Location: LABCELL_X18_Y65_N39
\TheRxFsk|Bandpasses:4:Bandpass0|Sample[-3]~12\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-3]~12_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a12~portbdataout\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ ) ) # ( 
-- \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a12~portbdataout\ & ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-3]~q\ ) ) ) # ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a12~portbdataout\ & ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-3]~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111000011110000111100000000000000001111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-3]~q\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a12~portbdataout\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-3]~12_combout\);

-- Location: FF_X16_Y63_N35
\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	asdata => \TheI2sToPar|D\(13),
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-2]~q\);

-- Location: LABCELL_X17_Y65_N33
\TheRxFsk|Bandpasses:4:Bandpass0|Sample[-2]~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-2]~13_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a13\ ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ 
-- & ( \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a13\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-2]~q\ ) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a13\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-2]~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111000000000000000000001111000011111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-2]~q\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a13\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-2]~13_combout\);

-- Location: LABCELL_X16_Y63_N15
\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-1]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-1]~feeder_combout\ = ( \TheI2sToPar|D\(14) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \TheI2sToPar|ALT_INV_D\(14),
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-1]~feeder_combout\);

-- Location: FF_X16_Y63_N16
\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-1]~feeder_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-1]~q\);

-- Location: LABCELL_X19_Y63_N12
\TheRxFsk|Bandpasses:4:Bandpass0|Sample[-1]~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-1]~14_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a14\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-1]~q\ ) ) # ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a14\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-1]~q\ & ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ ) ) ) # ( 
-- \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a14\ & ( !\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-1]~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000011110000111111110000111100001111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a14\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-1]~q\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|Sample[-1]~14_combout\);

-- Location: FF_X13_Y63_N37
\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[0]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	asdata => \TheI2sToPar|D\(15),
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[0]~DUPLICATE_q\);

-- Location: MLABCELL_X15_Y65_N51
\TheRxFsk|Bandpasses:4:Bandpass0|Sample[0]~15\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Sample[0]~15_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[0]~DUPLICATE_q\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a15\ ) ) # ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[0]~DUPLICATE_q\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a15\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ ) ) ) # ( 
-- \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[0]~DUPLICATE_q\ & ( !\TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a15\ & ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000001111000011111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[0]~DUPLICATE_q\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a15\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|Sample[0]~15_combout\);

-- Location: DSP_X20_Y65_N0
\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8\ : cyclonev_mac
-- pragma translate_off
GENERIC MAP (
	accumulate_clock => "none",
	ax_clock => "none",
	ax_width => 18,
	ay_scan_in_clock => "none",
	ay_scan_in_width => 19,
	ay_use_scan_in => "false",
	az_clock => "none",
	bx_clock => "none",
	by_clock => "none",
	by_use_scan_in => "false",
	bz_clock => "none",
	coef_a_0 => 0,
	coef_a_1 => 0,
	coef_a_2 => 0,
	coef_a_3 => 0,
	coef_a_4 => 0,
	coef_a_5 => 0,
	coef_a_6 => 0,
	coef_a_7 => 0,
	coef_b_0 => 0,
	coef_b_1 => 0,
	coef_b_2 => 0,
	coef_b_3 => 0,
	coef_b_4 => 0,
	coef_b_5 => 0,
	coef_b_6 => 0,
	coef_b_7 => 0,
	coef_sel_a_clock => "none",
	coef_sel_b_clock => "none",
	delay_scan_out_ay => "false",
	delay_scan_out_by => "false",
	enable_double_accum => "false",
	load_const_clock => "none",
	load_const_value => 0,
	mode_sub_location => 0,
	negate_clock => "none",
	operand_source_max => "input",
	operand_source_may => "input",
	operand_source_mbx => "input",
	operand_source_mby => "input",
	operation_mode => "m18x18_full",
	output_clock => "none",
	preadder_subtract_a => "false",
	preadder_subtract_b => "false",
	result_a_width => 64,
	signed_max => "true",
	signed_may => "true",
	signed_mbx => "false",
	signed_mby => "false",
	sub_clock => "none",
	use_chainadder => "false")
-- pragma translate_on
PORT MAP (
	sub => GND,
	negate => GND,
	ax => \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_AX_bus\,
	ay => \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_AY_bus\,
	resulta => \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_RESULTA_bus\);

-- Location: LABCELL_X18_Y65_N18
\TheRxFsk|Bandpasses:4:Bandpass0|vAdd~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|vAdd~2_combout\ = ( !\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~21\ & ( !\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~8_resulta\ & ( (!\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~12\ & (!\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~10\ & 
-- !\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~11\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1000000010000000000000000000000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~12\,
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~10\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~11\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~21\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~8_resulta\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|vAdd~2_combout\);

-- Location: MLABCELL_X21_Y65_N6
\TheRxFsk|Bandpasses:4:Bandpass0|vAdd~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|vAdd~1_combout\ = ( !\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~17\ & ( !\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~9\ & ( (!\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~14\ & (!\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~16\ & 
-- (!\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~15\ & !\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~18\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1000000000000000000000000000000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~14\,
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~16\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~15\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~18\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~17\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~9\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|vAdd~1_combout\);

-- Location: LABCELL_X19_Y65_N54
\TheRxFsk|Bandpasses:4:Bandpass0|vAdd~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|vAdd~0_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~13\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|vAdd~1_combout\ ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~13\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|vAdd~1_combout\ & 
-- ( (((!\TheRxFsk|Bandpasses:4:Bandpass0|vAdd~2_combout\) # (\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~22\)) # (\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~20\)) # (\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~19\) ) ) ) # ( \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~13\ & ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass0|vAdd~1_combout\ ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~13\ & ( !\TheRxFsk|Bandpasses:4:Bandpass0|vAdd~1_combout\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111111111111111111111111111111111111011111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~19\,
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~20\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~22\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_vAdd~2_combout\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~13\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_vAdd~1_combout\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|vAdd~0_combout\);

-- Location: LABCELL_X19_Y65_N0
\TheRxFsk|Bandpasses:4:Bandpass0|Add3~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add3~13_sumout\ = SUM(( (\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~39\ & \TheRxFsk|Bandpasses:4:Bandpass0|vAdd~0_combout\) ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~23\ ) + ( !VCC ))
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add3~14\ = CARRY(( (\TheRxFsk|Bandpasses:4:Bandpass0|Mult0~39\ & \TheRxFsk|Bandpasses:4:Bandpass0|vAdd~0_combout\) ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~23\ ) + ( !VCC ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111110000000000000000000000000000001100000011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~39\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_vAdd~0_combout\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~23\,
	cin => GND,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~13_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~14\);

-- Location: LABCELL_X19_Y65_N3
\TheRxFsk|Bandpasses:4:Bandpass0|Add3~17\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add3~17_sumout\ = SUM(( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~24\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add3~14\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add3~18\ = CARRY(( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~24\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add3~14\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~24\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~14\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~17_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~18\);

-- Location: LABCELL_X19_Y65_N6
\TheRxFsk|Bandpasses:4:Bandpass0|Add3~21\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add3~21_sumout\ = SUM(( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~25\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add3~18\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add3~22\ = CARRY(( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~25\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add3~18\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~25\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~18\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~21_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~22\);

-- Location: LABCELL_X19_Y65_N9
\TheRxFsk|Bandpasses:4:Bandpass0|Add3~25\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add3~25_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~26\ ) + ( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add3~22\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add3~26\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~26\ ) + ( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add3~22\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~26\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~22\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~25_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~26\);

-- Location: LABCELL_X19_Y65_N12
\TheRxFsk|Bandpasses:4:Bandpass0|Add3~29\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add3~29_sumout\ = SUM(( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~27\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add3~26\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add3~30\ = CARRY(( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~27\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add3~26\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~27\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~26\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~29_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~30\);

-- Location: LABCELL_X19_Y65_N15
\TheRxFsk|Bandpasses:4:Bandpass0|Add3~33\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add3~33_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~28\ ) + ( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add3~30\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add3~34\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~28\ ) + ( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add3~30\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~28\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~30\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~33_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~34\);

-- Location: LABCELL_X19_Y65_N18
\TheRxFsk|Bandpasses:4:Bandpass0|Add3~37\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add3~37_sumout\ = SUM(( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~29\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add3~34\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add3~38\ = CARRY(( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~29\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add3~34\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~29\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~34\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~37_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~38\);

-- Location: LABCELL_X19_Y65_N21
\TheRxFsk|Bandpasses:4:Bandpass0|Add3~41\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add3~41_sumout\ = SUM(( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~30\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add3~38\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add3~42\ = CARRY(( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~30\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add3~38\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~30\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~38\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~41_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~42\);

-- Location: LABCELL_X19_Y65_N24
\TheRxFsk|Bandpasses:4:Bandpass0|Add3~45\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add3~45_sumout\ = SUM(( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~31\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add3~42\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add3~46\ = CARRY(( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~31\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add3~42\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~31\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~42\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~45_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~46\);

-- Location: LABCELL_X19_Y65_N27
\TheRxFsk|Bandpasses:4:Bandpass0|Add3~49\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add3~49_sumout\ = SUM(( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~32\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add3~46\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add3~50\ = CARRY(( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~32\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add3~46\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~32\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~46\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~49_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~50\);

-- Location: LABCELL_X19_Y65_N30
\TheRxFsk|Bandpasses:4:Bandpass0|Add3~53\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add3~53_sumout\ = SUM(( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~33\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add3~50\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add3~54\ = CARRY(( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~33\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add3~50\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~33\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~50\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~53_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~54\);

-- Location: LABCELL_X19_Y65_N33
\TheRxFsk|Bandpasses:4:Bandpass0|Add3~57\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add3~57_sumout\ = SUM(( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~34\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add3~54\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add3~58\ = CARRY(( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~34\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add3~54\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~34\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~54\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~57_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~58\);

-- Location: LABCELL_X19_Y65_N36
\TheRxFsk|Bandpasses:4:Bandpass0|Add3~61\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add3~61_sumout\ = SUM(( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~35\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add3~58\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add3~62\ = CARRY(( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~35\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add3~58\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~35\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~58\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~61_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~62\);

-- Location: LABCELL_X19_Y65_N39
\TheRxFsk|Bandpasses:4:Bandpass0|Add3~65\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add3~65_sumout\ = SUM(( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~36\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add3~62\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add3~66\ = CARRY(( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~36\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add3~62\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000101010101010101000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~36\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~62\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~65_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~66\);

-- Location: LABCELL_X19_Y65_N42
\TheRxFsk|Bandpasses:4:Bandpass0|Add3~69\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add3~69_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~37\ ) + ( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add3~66\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add3~70\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~37\ ) + ( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add3~66\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~37\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~66\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~69_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~70\);

-- Location: LABCELL_X19_Y65_N45
\TheRxFsk|Bandpasses:4:Bandpass0|Add3~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add3~9_sumout\ = SUM(( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~38\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add3~70\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add3~10\ = CARRY(( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~38\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add3~70\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000101010101010101000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~38\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~70\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~9_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~10\);

-- Location: LABCELL_X19_Y65_N48
\TheRxFsk|Bandpasses:4:Bandpass0|Add3~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add3~5_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~39\ ) + ( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add3~10\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add3~6\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~39\ ) + ( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add3~10\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~39\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~10\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~5_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~6\);

-- Location: LABCELL_X19_Y65_N51
\TheRxFsk|Bandpasses:4:Bandpass0|Add3~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add3~1_sumout\ = SUM(( VCC ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Mult0~39\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add3~6\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000001111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Mult0~39\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~6\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~1_sumout\);

-- Location: LABCELL_X22_Y65_N54
\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[0]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[0]~0_combout\ = ( !\TheRxFsk|Bandpasses:4:Bandpass0|Add3~1_sumout\ )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111111111111111111111111111100000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add3~1_sumout\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[0]~0_combout\);

-- Location: FF_X22_Y65_N56
\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[0]~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed\(0));

-- Location: FF_X19_Y65_N46
\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_NEW_REG76\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~9_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM77\);

-- Location: FF_X19_Y65_N44
\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-1]_NEW_REG98\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~69_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-1]_OTERM99\);

-- Location: FF_X19_Y65_N49
\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_NEW_REG74\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~5_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM75\);

-- Location: FF_X19_Y65_N53
\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_NEW_REG72\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~1_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM73\);

-- Location: LABCELL_X23_Y65_N0
\TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-1]~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-1]~14_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM73\ & ( ((\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM75\) # 
-- (\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-1]_OTERM99\)) # (\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM77\) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM73\ & ( 
-- (\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM77\ & (\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-1]_OTERM99\ & \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM75\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000011000000000000001100111111111111110011111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM77\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-1]_OTERM99\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM75\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM73\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-1]~14_combout\);

-- Location: FF_X19_Y65_N40
\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-2]_NEW_REG104\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~65_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-2]_OTERM105\);

-- Location: MLABCELL_X21_Y65_N51
\TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-2]~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-2]~13_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-2]_OTERM105\ & ( ((\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM77\ & 
-- \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM75\)) # (\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM73\) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-2]_OTERM105\ & ( 
-- (\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM73\ & ((\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM75\) # (\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM77\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001001100010011000100110001001100110111001101110011011100110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM77\,
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM73\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM75\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-2]_OTERM105\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-2]~13_combout\);

-- Location: FF_X19_Y65_N37
\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-3]_NEW_REG110\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~61_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-3]_OTERM111\);

-- Location: MLABCELL_X21_Y65_N48
\TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-3]~12\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-3]~12_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-3]_OTERM111\ & ( ((\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM77\ & 
-- \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM75\)) # (\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM73\) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-3]_OTERM111\ & ( 
-- (\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM73\ & ((\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM75\) # (\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM77\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000100110011000100010011001100110011011101110011001101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM77\,
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM73\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM75\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-3]_OTERM111\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-3]~12_combout\);

-- Location: FF_X19_Y65_N34
\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-4]_NEW_REG116\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~57_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-4]_OTERM117\);

-- Location: MLABCELL_X21_Y65_N33
\TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-4]~11\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-4]~11_combout\ = (!\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM77\ & (\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM73\ & 
-- ((\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM75\) # (\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-4]_OTERM117\)))) # (\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM77\ & 
-- (((\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-4]_OTERM117\ & \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM75\)) # (\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM73\)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001001100110111000100110011011100010011001101110001001100110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM77\,
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM73\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-4]_OTERM117\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM75\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-4]~11_combout\);

-- Location: FF_X19_Y65_N31
\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-5]_NEW_REG122\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~53_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-5]_OTERM123\);

-- Location: MLABCELL_X21_Y65_N30
\TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-5]~10\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-5]~10_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-5]_OTERM123\ & ( ((\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM77\ & 
-- \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM75\)) # (\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM73\) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-5]_OTERM123\ & ( 
-- (\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM73\ & ((\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM75\) # (\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM77\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000100110011000100010011001100110011011101110011001101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM77\,
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM73\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM75\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-5]_OTERM123\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-5]~10_combout\);

-- Location: FF_X19_Y65_N28
\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-6]_NEW_REG128\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~49_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-6]_OTERM129\);

-- Location: MLABCELL_X21_Y65_N39
\TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-6]~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-6]~9_combout\ = (!\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM77\ & (\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM73\ & 
-- ((\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM75\) # (\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-6]_OTERM129\)))) # (\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM77\ & 
-- (((\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-6]_OTERM129\ & \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM75\)) # (\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM73\)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001001100110111000100110011011100010011001101110001001100110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM77\,
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM73\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-6]_OTERM129\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM75\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-6]~9_combout\);

-- Location: FF_X19_Y65_N25
\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-7]_NEW_REG134\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~45_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-7]_OTERM135\);

-- Location: MLABCELL_X21_Y65_N36
\TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-7]~8\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-7]~8_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-7]_OTERM135\ & ( ((\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM77\ & 
-- \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM75\)) # (\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM73\) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-7]_OTERM135\ & ( 
-- (\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM73\ & ((\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM75\) # (\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM77\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000100110011000100010011001100110011011101110011001101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM77\,
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM73\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM75\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-7]_OTERM135\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-7]~8_combout\);

-- Location: FF_X19_Y65_N22
\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-8]_NEW_REG140\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~41_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-8]_OTERM141\);

-- Location: MLABCELL_X21_Y65_N21
\TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-8]~7\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-8]~7_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM75\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-8]_OTERM141\ & ( 
-- (\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM73\) # (\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM77\) ) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM75\ & ( 
-- \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-8]_OTERM141\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM73\ ) ) ) # ( \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM75\ & ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-8]_OTERM141\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM73\ ) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM75\ & ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-8]_OTERM141\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM77\ & \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM73\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100000101000011110000111100001111000011110101111101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM77\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM73\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM75\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-8]_OTERM141\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-8]~7_combout\);

-- Location: FF_X19_Y65_N19
\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-9]_NEW_REG146\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~37_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-9]_OTERM147\);

-- Location: MLABCELL_X21_Y65_N0
\TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-9]~6\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-9]~6_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM75\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-9]_OTERM147\ & ( 
-- (\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM77\) # (\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM73\) ) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM75\ & ( 
-- \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-9]_OTERM147\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM73\ ) ) ) # ( \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM75\ & ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-9]_OTERM147\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM73\ ) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM75\ & ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-9]_OTERM147\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM73\ & \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM77\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100000011001100110011001100110011001100110011111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM73\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM77\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM75\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-9]_OTERM147\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-9]~6_combout\);

-- Location: FF_X19_Y65_N16
\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-10]_NEW_REG152\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~33_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-10]_OTERM153\);

-- Location: MLABCELL_X21_Y65_N45
\TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-10]~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-10]~5_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-10]_OTERM153\ & ( ((\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM77\ & 
-- \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM75\)) # (\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM73\) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-10]_OTERM153\ & ( 
-- (\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM73\ & ((\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM75\) # (\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM77\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000011100000111000111110001111100000111000001110001111100011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM77\,
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM75\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM73\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-10]_OTERM153\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-10]~5_combout\);

-- Location: FF_X19_Y65_N13
\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-11]_NEW_REG158\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~29_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-11]_OTERM159\);

-- Location: MLABCELL_X21_Y65_N12
\TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-11]~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-11]~4_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM75\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-11]_OTERM159\ & ( 
-- (\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM77\) # (\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM73\) ) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM75\ & ( 
-- \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-11]_OTERM159\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM73\ ) ) ) # ( \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM75\ & ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-11]_OTERM159\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM73\ ) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM75\ & ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-11]_OTERM159\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM73\ & \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM77\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100000011001100110011001100110011001100110011111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM73\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM77\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM75\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-11]_OTERM159\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-11]~4_combout\);

-- Location: FF_X19_Y65_N10
\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-12]_NEW_REG164\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~25_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-12]_OTERM165\);

-- Location: MLABCELL_X21_Y65_N57
\TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-12]~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-12]~3_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-12]_OTERM165\ & ( ((\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM77\ & 
-- \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM75\)) # (\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM73\) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-12]_OTERM165\ & ( 
-- (\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM73\ & ((\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM75\) # (\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM77\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000011100000111000001110000011100011111000111110001111100011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM77\,
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM75\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM73\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-12]_OTERM165\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-12]~3_combout\);

-- Location: FF_X19_Y65_N8
\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-13]_NEW_REG170\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~21_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-13]_OTERM171\);

-- Location: MLABCELL_X21_Y65_N24
\TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-13]~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-13]~2_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM73\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-13]_OTERM171\ ) ) # ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM73\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-13]_OTERM171\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM77\ & 
-- \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM75\) ) ) ) # ( \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM73\ & ( !\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-13]_OTERM171\ & ( 
-- (\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM75\) # (\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM77\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000011111111111100000000000011111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM77\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM75\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM73\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-13]_OTERM171\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-13]~2_combout\);

-- Location: FF_X19_Y65_N5
\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-14]_NEW_REG176\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~17_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-14]_OTERM177\);

-- Location: LABCELL_X18_Y65_N12
\TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-14]~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-14]~1_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM75\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM73\ ) ) # ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM75\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM73\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM77\) # 
-- (\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-14]_OTERM177\) ) ) ) # ( \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM75\ & ( !\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM73\ & ( 
-- (\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-14]_OTERM177\ & \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM77\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000001010000010101011111010111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-14]_OTERM177\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM77\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM75\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM73\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-14]~1_combout\);

-- Location: FF_X19_Y65_N1
\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_NEW_REG78\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|Add3~13_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM79\);

-- Location: LABCELL_X23_Y65_N9
\TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-15]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-15]~0_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM79\ & ( ((\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM75\ & 
-- \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM77\)) # (\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM73\) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM79\ & ( 
-- (\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM73\ & ((\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM77\) # (\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed[-15]_OTERM75\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010101010101000001010101010101010101010111110101010101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM73\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM75\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM77\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM79\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-15]~0_combout\);

-- Location: LABCELL_X22_Y65_N45
\TheRxFsk|Bandpasses:4:Bandpass0|Add4~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add4~5_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass0|Sum\(0) ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed\(0) ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add4~66\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add4~6\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass0|Sum\(0) ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed\(0) ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add4~66\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000101010101010101000000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed\(0),
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum\(0),
	cin => \TheRxFsk|Bandpasses:4:Bandpass0|Add4~66\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass0|Add4~5_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass0|Add4~6\);

-- Location: LABCELL_X23_Y65_N6
\TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-15]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-15]~0_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|Add4~5_sumout\ & ( (!\TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-15]~0_combout\ $ (!\TheRxFsk|Bandpasses:4:Bandpass0|Sum[-15]~q\)) # 
-- (\TheRxFsk|Bandpasses:4:Bandpass0|Add4~1_sumout\) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|Add4~1_sumout\ & (!\TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-15]~0_combout\ $ 
-- (!\TheRxFsk|Bandpasses:4:Bandpass0|Sum[-15]~q\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100110000000000110011000000111111111100110011111111110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~1_sumout\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResult[-15]~0_combout\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-15]~q\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~5_sumout\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-15]~0_combout\);

-- Location: LABCELL_X16_Y61_N42
\TheRxFsk|Bandpasses:4:Bandpass0|Selector2~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Selector2~0_combout\ = ( \TheRxFsk|Bandpasses:11:Bandpass1|Equal1~1_combout\ & ( ((!\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~0_combout\ & \TheRxFsk|Bandpasses:4:Bandpass0|R.SumState.SumSelect~q\)) # 
-- (\TheRxFsk|Bandpasses:4:Bandpass0|R.SumState.SumEnable~q\) ) ) # ( !\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~1_combout\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|R.SumState.SumSelect~q\) # (\TheRxFsk|Bandpasses:4:Bandpass0|R.SumState.SumEnable~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111111111111000011111111111100001111101011110000111110101111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:11:Bandpass1|ALT_INV_Equal1~0_combout\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.SumState.SumEnable~q\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.SumState.SumSelect~q\,
	dataf => \TheRxFsk|Bandpasses:11:Bandpass1|ALT_INV_Equal1~1_combout\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|Selector2~0_combout\);

-- Location: FF_X16_Y61_N44
\TheRxFsk|Bandpasses:4:Bandpass0|R.SumState.SumSelect\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|Selector2~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|R.SumState.SumSelect~q\);

-- Location: LABCELL_X16_Y61_N45
\TheRxFsk|Bandpasses:4:Bandpass0|Selector3~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Selector3~0_combout\ = ( \TheRxFsk|Bandpasses:11:Bandpass1|Equal1~1_combout\ & ( (\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~0_combout\ & \TheRxFsk|Bandpasses:4:Bandpass0|R.SumState.SumSelect~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000101000001010000010100000101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:11:Bandpass1|ALT_INV_Equal1~0_combout\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.SumState.SumSelect~q\,
	dataf => \TheRxFsk|Bandpasses:11:Bandpass1|ALT_INV_Equal1~1_combout\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|Selector3~0_combout\);

-- Location: FF_X16_Y61_N47
\TheRxFsk|Bandpasses:4:Bandpass0|R.SumState.SumWait1\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|Selector3~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|R.SumState.SumWait1~q\);

-- Location: FF_X16_Y61_N41
\TheRxFsk|Bandpasses:4:Bandpass0|R.SumState.SumWait2\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	asdata => \TheRxFsk|Bandpasses:4:Bandpass0|R.SumState.SumWait1~q\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|R.SumState.SumWait2~q\);

-- Location: FF_X16_Y61_N50
\TheRxFsk|Bandpasses:4:Bandpass0|R.SumState.SumValid\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	asdata => \TheRxFsk|Bandpasses:4:Bandpass0|R.SumState.SumWait2~q\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|R.SumState.SumValid~q\);

-- Location: LABCELL_X16_Y61_N0
\TheRxFsk|Bandpasses:4:Bandpass0|Selector0~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Selector0~0_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|R.SumState.Idle~q\ & ( \TheI2sToPar|ValL~q\ & ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.SumState.SumValid~q\ ) ) ) # ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass0|R.SumState.Idle~q\ & ( \TheI2sToPar|ValL~q\ & ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.SumState.SumValid~q\ ) ) ) # ( \TheRxFsk|Bandpasses:4:Bandpass0|R.SumState.Idle~q\ & ( !\TheI2sToPar|ValL~q\ & ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass0|R.SumState.SumValid~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000011110000111100001111000011110000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.SumState.SumValid~q\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.SumState.Idle~q\,
	dataf => \TheI2sToPar|ALT_INV_ValL~q\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|Selector0~0_combout\);

-- Location: FF_X16_Y61_N2
\TheRxFsk|Bandpasses:4:Bandpass0|R.SumState.Idle\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|Selector0~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|R.SumState.Idle~q\);

-- Location: LABCELL_X16_Y61_N33
\TheRxFsk|Bandpasses:4:Bandpass0|Selector1~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Selector1~0_combout\ = ( \TheI2sToPar|ValL~q\ & ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.SumState.Idle~q\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000010101010101010101010101010101010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.SumState.Idle~q\,
	dataf => \TheI2sToPar|ALT_INV_ValL~q\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|Selector1~0_combout\);

-- Location: FF_X16_Y61_N35
\TheRxFsk|Bandpasses:4:Bandpass0|R.SumState.SumEnable\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|Selector1~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|R.SumState.SumEnable~q\);

-- Location: LABCELL_X16_Y61_N12
\TheRxFsk|Bandpasses:4:Bandpass0|Selector6~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Selector6~0_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|R.SelSumUp~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|R.SumState.SumWait2~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|R.SumState.SumEnable~q\ ) ) ) # ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass0|R.SelSumUp~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|R.SumState.SumWait2~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|R.SumState.SumEnable~q\ ) ) ) # ( \TheRxFsk|Bandpasses:4:Bandpass0|R.SelSumUp~q\ & ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass0|R.SumState.SumWait2~q\ ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.SelSumUp~q\ & ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.SumState.SumWait2~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|R.SumState.SumEnable~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111111111111111111100001111000011110000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.SumState.SumEnable~q\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.SelSumUp~q\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.SumState.SumWait2~q\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|Selector6~0_combout\);

-- Location: FF_X16_Y61_N13
\TheRxFsk|Bandpasses:4:Bandpass0|R.SelSumUp\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|Selector6~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|R.SelSumUp~q\);

-- Location: LABCELL_X16_Y61_N6
\TheRxFsk|Bandpasses:4:Bandpass0|Selector7~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Selector7~0_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|R.EnableSumUp~q\ & ( \TheI2sToPar|ValL~q\ & ( (!\TheRxFsk|Bandpasses:4:Bandpass0|R.SumState.Idle~q\) # (!\TheRxFsk|Bandpasses:4:Bandpass0|R.SumState.SumWait2~q\) ) 
-- ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.EnableSumUp~q\ & ( \TheI2sToPar|ValL~q\ & ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.SumState.Idle~q\ ) ) ) # ( \TheRxFsk|Bandpasses:4:Bandpass0|R.EnableSumUp~q\ & ( !\TheI2sToPar|ValL~q\ & ( 
-- (!\TheRxFsk|Bandpasses:4:Bandpass0|R.SumState.Idle~q\) # (!\TheRxFsk|Bandpasses:4:Bandpass0|R.SumState.SumWait2~q\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111000011110000111100001111111111110000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.SumState.Idle~q\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.SumState.SumWait2~q\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.EnableSumUp~q\,
	dataf => \TheI2sToPar|ALT_INV_ValL~q\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|Selector7~0_combout\);

-- Location: FF_X16_Y61_N7
\TheRxFsk|Bandpasses:4:Bandpass0|R.EnableSumUp\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|Selector7~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|R.EnableSumUp~q\);

-- Location: FF_X23_Y65_N7
\TheRxFsk|Bandpasses:4:Bandpass0|Sum[-15]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-15]~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:4:Bandpass0|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-15]~q\);

-- Location: LABCELL_X22_Y65_N0
\TheRxFsk|Bandpasses:4:Bandpass0|Add4~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add4~10\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-15]~0_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-15]~q\ ) + ( !VCC ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000110011001100110000000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-15]~q\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResult[-15]~0_combout\,
	cin => GND,
	cout => \TheRxFsk|Bandpasses:4:Bandpass0|Add4~10\);

-- Location: LABCELL_X22_Y65_N3
\TheRxFsk|Bandpasses:4:Bandpass0|Add4~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add4~13_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-14]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-14]~1_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add4~10\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add4~14\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-14]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-14]~1_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add4~10\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-14]~q\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResult[-14]~1_combout\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass0|Add4~10\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass0|Add4~13_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass0|Add4~14\);

-- Location: LABCELL_X23_Y65_N15
\TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-14]~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-14]~1_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|Add4~13_sumout\) # (\TheRxFsk|Bandpasses:4:Bandpass0|Add4~1_sumout\) ) ) # ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass0|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|Add4~1_sumout\ & \TheRxFsk|Bandpasses:4:Bandpass0|Add4~13_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100000011000000110000001100111111001111110011111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~1_sumout\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~13_sumout\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~5_sumout\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-14]~1_combout\);

-- Location: FF_X23_Y65_N16
\TheRxFsk|Bandpasses:4:Bandpass0|Sum[-14]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-14]~1_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:4:Bandpass0|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-14]~q\);

-- Location: LABCELL_X22_Y65_N6
\TheRxFsk|Bandpasses:4:Bandpass0|Add4~17\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add4~17_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-13]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-13]~2_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add4~14\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add4~18\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-13]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-13]~2_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add4~14\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000110011001100110000000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResult[-13]~2_combout\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-13]~q\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass0|Add4~14\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass0|Add4~17_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass0|Add4~18\);

-- Location: LABCELL_X23_Y65_N30
\TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-13]~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-13]~2_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|Add4~17_sumout\) # (\TheRxFsk|Bandpasses:4:Bandpass0|Add4~1_sumout\) ) ) # ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass0|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|Add4~1_sumout\ & \TheRxFsk|Bandpasses:4:Bandpass0|Add4~17_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100000011000000110000001100111111001111110011111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~1_sumout\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~17_sumout\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~5_sumout\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-13]~2_combout\);

-- Location: FF_X23_Y65_N32
\TheRxFsk|Bandpasses:4:Bandpass0|Sum[-13]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-13]~2_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:4:Bandpass0|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-13]~q\);

-- Location: LABCELL_X22_Y65_N9
\TheRxFsk|Bandpasses:4:Bandpass0|Add4~21\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add4~21_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-12]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-12]~3_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add4~18\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add4~22\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-12]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-12]~3_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add4~18\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-12]~q\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResult[-12]~3_combout\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass0|Add4~18\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass0|Add4~21_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass0|Add4~22\);

-- Location: LABCELL_X23_Y65_N33
\TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-12]~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-12]~3_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|Add4~21_sumout\) # (\TheRxFsk|Bandpasses:4:Bandpass0|Add4~1_sumout\) ) ) # ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass0|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|Add4~1_sumout\ & \TheRxFsk|Bandpasses:4:Bandpass0|Add4~21_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000110011000000000011001100110011111111110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~1_sumout\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~21_sumout\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~5_sumout\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-12]~3_combout\);

-- Location: FF_X23_Y65_N34
\TheRxFsk|Bandpasses:4:Bandpass0|Sum[-12]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-12]~3_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:4:Bandpass0|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-12]~q\);

-- Location: LABCELL_X22_Y65_N12
\TheRxFsk|Bandpasses:4:Bandpass0|Add4~25\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add4~25_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-11]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-11]~4_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add4~22\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add4~26\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-11]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-11]~4_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add4~22\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-11]~q\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResult[-11]~4_combout\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass0|Add4~22\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass0|Add4~25_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass0|Add4~26\);

-- Location: LABCELL_X23_Y65_N24
\TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-11]~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-11]~4_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|Add4~25_sumout\) # (\TheRxFsk|Bandpasses:4:Bandpass0|Add4~1_sumout\) ) ) # ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass0|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|Add4~1_sumout\ & \TheRxFsk|Bandpasses:4:Bandpass0|Add4~25_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100000011000000110000001100111111001111110011111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~1_sumout\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~25_sumout\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~5_sumout\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-11]~4_combout\);

-- Location: FF_X23_Y65_N25
\TheRxFsk|Bandpasses:4:Bandpass0|Sum[-11]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-11]~4_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:4:Bandpass0|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-11]~q\);

-- Location: LABCELL_X22_Y65_N15
\TheRxFsk|Bandpasses:4:Bandpass0|Add4~29\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add4~29_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-10]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-10]~5_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add4~26\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add4~30\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-10]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-10]~5_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add4~26\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111110000000000000000000000000101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-10]~q\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResult[-10]~5_combout\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass0|Add4~26\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass0|Add4~29_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass0|Add4~30\);

-- Location: LABCELL_X23_Y65_N27
\TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-10]~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-10]~5_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|Add4~29_sumout\) # (\TheRxFsk|Bandpasses:4:Bandpass0|Add4~1_sumout\) ) ) # ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass0|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|Add4~1_sumout\ & \TheRxFsk|Bandpasses:4:Bandpass0|Add4~29_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100000011000000110000001100111111001111110011111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~1_sumout\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~29_sumout\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~5_sumout\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-10]~5_combout\);

-- Location: FF_X23_Y65_N29
\TheRxFsk|Bandpasses:4:Bandpass0|Sum[-10]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-10]~5_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:4:Bandpass0|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-10]~q\);

-- Location: LABCELL_X22_Y65_N18
\TheRxFsk|Bandpasses:4:Bandpass0|Add4~33\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add4~33_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-9]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-9]~6_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add4~30\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add4~34\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-9]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-9]~6_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add4~30\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000110011001100110000000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResult[-9]~6_combout\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-9]~q\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass0|Add4~30\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass0|Add4~33_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass0|Add4~34\);

-- Location: LABCELL_X23_Y65_N54
\TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-9]~6\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-9]~6_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|Add4~33_sumout\) # (\TheRxFsk|Bandpasses:4:Bandpass0|Add4~1_sumout\) ) ) # ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass0|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|Add4~1_sumout\ & \TheRxFsk|Bandpasses:4:Bandpass0|Add4~33_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100000011000000110000001100111111001111110011111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~1_sumout\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~33_sumout\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~5_sumout\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-9]~6_combout\);

-- Location: FF_X23_Y65_N56
\TheRxFsk|Bandpasses:4:Bandpass0|Sum[-9]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-9]~6_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:4:Bandpass0|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-9]~q\);

-- Location: LABCELL_X22_Y65_N21
\TheRxFsk|Bandpasses:4:Bandpass0|Add4~37\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add4~37_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-8]~7_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-8]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add4~34\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add4~38\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-8]~7_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-8]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add4~34\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000101010101010101000000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-8]~q\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResult[-8]~7_combout\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass0|Add4~34\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass0|Add4~37_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass0|Add4~38\);

-- Location: LABCELL_X23_Y65_N57
\TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-8]~7\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-8]~7_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|Add4~37_sumout\) # (\TheRxFsk|Bandpasses:4:Bandpass0|Add4~1_sumout\) ) ) # ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass0|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|Add4~1_sumout\ & \TheRxFsk|Bandpasses:4:Bandpass0|Add4~37_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000110011000000000011001100110011111111110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~1_sumout\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~37_sumout\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~5_sumout\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-8]~7_combout\);

-- Location: FF_X23_Y65_N58
\TheRxFsk|Bandpasses:4:Bandpass0|Sum[-8]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-8]~7_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:4:Bandpass0|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-8]~q\);

-- Location: LABCELL_X22_Y65_N24
\TheRxFsk|Bandpasses:4:Bandpass0|Add4~41\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add4~41_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-7]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-7]~8_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add4~38\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add4~42\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-7]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-7]~8_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add4~38\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111110000000000000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-7]~q\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResult[-7]~8_combout\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass0|Add4~38\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass0|Add4~41_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass0|Add4~42\);

-- Location: LABCELL_X23_Y65_N3
\TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-7]~8\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-7]~8_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|Add4~1_sumout\) # (\TheRxFsk|Bandpasses:4:Bandpass0|Add4~41_sumout\) ) ) # ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass0|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|Add4~41_sumout\ & \TheRxFsk|Bandpasses:4:Bandpass0|Add4~1_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000001111000000000000111100001111111111110000111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~41_sumout\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~1_sumout\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~5_sumout\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-7]~8_combout\);

-- Location: FF_X23_Y65_N5
\TheRxFsk|Bandpasses:4:Bandpass0|Sum[-7]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-7]~8_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:4:Bandpass0|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-7]~q\);

-- Location: LABCELL_X22_Y65_N27
\TheRxFsk|Bandpasses:4:Bandpass0|Add4~45\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add4~45_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-6]~9_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-6]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add4~42\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add4~46\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-6]~9_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-6]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add4~42\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111110000000000000000000000000101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResult[-6]~9_combout\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-6]~q\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass0|Add4~42\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass0|Add4~45_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass0|Add4~46\);

-- Location: LABCELL_X23_Y65_N45
\TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-6]~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-6]~9_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|Add4~45_sumout\) # (\TheRxFsk|Bandpasses:4:Bandpass0|Add4~1_sumout\) ) ) # ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass0|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|Add4~1_sumout\ & \TheRxFsk|Bandpasses:4:Bandpass0|Add4~45_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000110011000000000011001100110011111111110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~1_sumout\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~45_sumout\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~5_sumout\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-6]~9_combout\);

-- Location: FF_X23_Y65_N47
\TheRxFsk|Bandpasses:4:Bandpass0|Sum[-6]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-6]~9_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:4:Bandpass0|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-6]~q\);

-- Location: LABCELL_X22_Y65_N30
\TheRxFsk|Bandpasses:4:Bandpass0|Add4~49\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add4~49_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-5]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-5]~10_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add4~46\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add4~50\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-5]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-5]~10_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add4~46\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResult[-5]~10_combout\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-5]~q\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass0|Add4~46\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass0|Add4~49_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass0|Add4~50\);

-- Location: LABCELL_X23_Y65_N36
\TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-5]~10\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-5]~10_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|Add4~49_sumout\) # (\TheRxFsk|Bandpasses:4:Bandpass0|Add4~1_sumout\) ) ) # ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass0|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|Add4~1_sumout\ & \TheRxFsk|Bandpasses:4:Bandpass0|Add4~49_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100000011000000110000001100111111001111110011111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~1_sumout\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~49_sumout\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~5_sumout\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-5]~10_combout\);

-- Location: FF_X23_Y65_N37
\TheRxFsk|Bandpasses:4:Bandpass0|Sum[-5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-5]~10_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:4:Bandpass0|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-5]~q\);

-- Location: LABCELL_X22_Y65_N33
\TheRxFsk|Bandpasses:4:Bandpass0|Add4~53\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add4~53_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-4]~11_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-4]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add4~50\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add4~54\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-4]~11_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-4]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add4~50\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111110000000000000000000000000011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResult[-4]~11_combout\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-4]~q\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass0|Add4~50\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass0|Add4~53_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass0|Add4~54\);

-- Location: LABCELL_X23_Y65_N39
\TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-4]~11\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-4]~11_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|Add4~53_sumout\) # (\TheRxFsk|Bandpasses:4:Bandpass0|Add4~1_sumout\) ) ) # ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass0|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|Add4~1_sumout\ & \TheRxFsk|Bandpasses:4:Bandpass0|Add4~53_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100000011000000110000001100111111001111110011111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~1_sumout\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~53_sumout\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~5_sumout\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-4]~11_combout\);

-- Location: FF_X23_Y65_N41
\TheRxFsk|Bandpasses:4:Bandpass0|Sum[-4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-4]~11_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:4:Bandpass0|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-4]~q\);

-- Location: LABCELL_X22_Y65_N36
\TheRxFsk|Bandpasses:4:Bandpass0|Add4~57\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add4~57_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-3]~12_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-3]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add4~54\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add4~58\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-3]~12_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-3]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add4~54\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000110011001100110000000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-3]~q\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResult[-3]~12_combout\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass0|Add4~54\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass0|Add4~57_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass0|Add4~58\);

-- Location: LABCELL_X23_Y65_N18
\TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-3]~12\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-3]~12_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|Add4~57_sumout\) # (\TheRxFsk|Bandpasses:4:Bandpass0|Add4~1_sumout\) ) ) # ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass0|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|Add4~1_sumout\ & \TheRxFsk|Bandpasses:4:Bandpass0|Add4~57_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100000011000000110000001100111111001111110011111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~1_sumout\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~57_sumout\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~5_sumout\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-3]~12_combout\);

-- Location: FF_X23_Y65_N20
\TheRxFsk|Bandpasses:4:Bandpass0|Sum[-3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-3]~12_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:4:Bandpass0|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-3]~q\);

-- Location: LABCELL_X22_Y65_N39
\TheRxFsk|Bandpasses:4:Bandpass0|Add4~61\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add4~61_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-2]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-2]~13_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add4~58\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add4~62\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-2]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-2]~13_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add4~58\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111110000000000000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-2]~q\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResult[-2]~13_combout\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass0|Add4~58\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass0|Add4~61_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass0|Add4~62\);

-- Location: LABCELL_X23_Y65_N21
\TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-2]~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-2]~13_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|Add4~1_sumout\) # (\TheRxFsk|Bandpasses:4:Bandpass0|Add4~61_sumout\) ) ) # ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass0|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|Add4~61_sumout\ & \TheRxFsk|Bandpasses:4:Bandpass0|Add4~1_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000100010001000100010001000101110111011101110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~61_sumout\,
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~1_sumout\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~5_sumout\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-2]~13_combout\);

-- Location: FF_X23_Y65_N22
\TheRxFsk|Bandpasses:4:Bandpass0|Sum[-2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-2]~13_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:4:Bandpass0|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-2]~q\);

-- Location: LABCELL_X22_Y65_N42
\TheRxFsk|Bandpasses:4:Bandpass0|Add4~65\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add4~65_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-1]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-1]~14_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add4~62\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add4~66\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-1]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|MultResult[-1]~14_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add4~62\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-1]~q\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResult[-1]~14_combout\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass0|Add4~62\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass0|Add4~65_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass0|Add4~66\);

-- Location: LABCELL_X23_Y65_N42
\TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-1]~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-1]~14_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|Add4~65_sumout\) # (\TheRxFsk|Bandpasses:4:Bandpass0|Add4~1_sumout\) ) ) # ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass0|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|Add4~1_sumout\ & \TheRxFsk|Bandpasses:4:Bandpass0|Add4~65_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000110011000000000011001100110011111111110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~1_sumout\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~65_sumout\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~5_sumout\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-1]~14_combout\);

-- Location: FF_X23_Y65_N44
\TheRxFsk|Bandpasses:4:Bandpass0|Sum[-1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|NextSum[-1]~14_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:4:Bandpass0|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-1]~q\);

-- Location: LABCELL_X22_Y65_N48
\TheRxFsk|Bandpasses:4:Bandpass0|Add4~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add4~1_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass0|Sum\(0) ) + ( !\TheRxFsk|Bandpasses:4:Bandpass0|MultResultDelayed\(0) ) + ( \TheRxFsk|Bandpasses:4:Bandpass0|Add4~6\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000011110000111100000000000000000011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum\(0),
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_MultResultDelayed\(0),
	cin => \TheRxFsk|Bandpasses:4:Bandpass0|Add4~6\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass0|Add4~1_sumout\);

-- Location: LABCELL_X23_Y65_N48
\TheRxFsk|Bandpasses:4:Bandpass0|Add4~1_wirecell\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass0|Add4~1_wirecell_combout\ = ( !\TheRxFsk|Bandpasses:4:Bandpass0|Add4~1_sumout\ )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111111111111000000000000000011111111111111110000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Add4~1_sumout\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass0|Add4~1_wirecell_combout\);

-- Location: FF_X23_Y65_N49
\TheRxFsk|Bandpasses:4:Bandpass0|Sum[0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass0|Add4~1_wirecell_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:4:Bandpass0|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|Sum\(0));

-- Location: M10K_X26_Y59_N0
\TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a4\ : cyclonev_ram_block
-- pragma translate_off
GENERIC MAP (
	mem_init4 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	mem_init3 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	mem_init2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001D00241003EAFFDF2FFFEC0010A0001BFFE0F000EE001DEFFFF6FFE1D0012500101FFDD8FFFDA0020A00033FFC22000E6003C3FFEE6FFC2B003430020CFFBC2FFEBB0040500050FFA41001E3005A0FFCCAFFB370046B00323FF9ACFFE90007F7FFF6FFF86C002E900778FFAA0FF93C0079B00448FF69BFFD5B00ADAFFF8CFF5A4004FC00A4",
	mem_init1 => "FFF869FF73500ACD0057BFF395FFD2100DADFFEA1FF1E30061E00C2DFF528FF51F00DFC006BBFEF9DFFDE701172FFCA7FEE250085100F17FF2E2FF4F80112000703FECB7FFEB60152CFFB9CFEB6100A9101113FEF9EFF2C0014330074BFE8E4FFF94018E2FF97CFE98F00DD901325FEC65FF27D017310068CFE51F0008801A9CFF74AFE7A900F220144BFEA3EFF23501A17006BDFE3640029501C62FF50BFE6AA0116201483FE830FF2F001BE8005D8FE2AA003B901C3DFF4C6FE69101391013C6FE63DFF4B901CAA003D8FE2E8005F001B30FF283FE862014AA0110BFE662FF59501C64002BDFE3170063501A3EFF24BFEA22014A900F4AFE79CFF78801A1F0",
	mem_init0 => "008CFE5310067D01765FF225FECD90138F00D7CFE9E2FF994018E4FFF4BFE833007C00149EFF213FEF910116100A9CFEB2CFFBB6015B7FFE03FEC20007F8011E2FF417FF25100F25008A7FEE72FFCE70119DFFDBBFEFFC0061F00D28FF52DFF51E00CE3006A1FF1ADFFE2100D95FFD7BFF3CD0053500A69FF74FFF8FC00AA40048CFF5DAFFF5B00A9BFFD48FF69B0043C007A0FF978FFAE90076C0026FFF8F7FFF90007ACFFE23FF96B00337004CAFFBA0FFCE30054100150FFA05000BB004C2FFE0CFFB430022B003E6FFCC3FFEE60032200033FFC0A000DA002D8FFF01FFD250011D001F6FFEDEFFFEE0010F0001BFFE0A000EC001F2FFFEAFFD410031D002",
	data_interleave_offset_in_bits => 1,
	data_interleave_width_in_bits => 1,
	init_file => "db/TbdRxFskBasic.ram1_DspFir_2df41c30.hdl.mif",
	init_file_layout => "port_a",
	logical_ram_name => "RxFsk:TheRxFsk|DspFir:\Bandpasses:4:Bandpass1|altsyncram:CoefMemory_rtl_0|altsyncram_2nd1:auto_generated|ALTSYNCRAM",
	operation_mode => "rom",
	port_a_address_clear => "none",
	port_a_address_width => 9,
	port_a_byte_enable_clock => "none",
	port_a_data_out_clear => "none",
	port_a_data_out_clock => "none",
	port_a_data_width => 20,
	port_a_first_address => 0,
	port_a_first_bit_number => 0,
	port_a_last_address => 511,
	port_a_logical_ram_depth => 258,
	port_a_logical_ram_width => 16,
	port_a_read_during_write_mode => "new_data_no_nbe_read",
	port_a_write_enable_clock => "none",
	port_b_address_width => 9,
	port_b_data_width => 20,
	ram_block_type => "M20K")
-- pragma translate_on
PORT MAP (
	portare => VCC,
	clk0 => \iClk~inputCLKENA0_outclk\,
	portaaddr => \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a4_PORTAADDR_bus\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	portadataout => \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a4_PORTADATAOUT_bus\);

-- Location: M10K_X14_Y62_N0
\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a4\ : cyclonev_ram_block
-- pragma translate_off
GENERIC MAP (
	mem_init4 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	mem_init3 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	mem_init2 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	mem_init1 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	mem_init0 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	data_interleave_offset_in_bits => 1,
	data_interleave_width_in_bits => 1,
	init_file => "db/TbdRxFskBasic.ram0_DspFir_2df41c30.hdl.mif",
	init_file_layout => "port_a",
	logical_ram_name => "RxFsk:TheRxFsk|DspFir:\Bandpasses:4:Bandpass1|altsyncram:SampleMemory_rtl_0|altsyncram_cbs1:auto_generated|ALTSYNCRAM",
	mixed_port_feed_through_mode => "old",
	operation_mode => "dual_port",
	port_a_address_clear => "none",
	port_a_address_width => 9,
	port_a_byte_enable_clock => "none",
	port_a_data_out_clear => "none",
	port_a_data_out_clock => "none",
	port_a_data_width => 20,
	port_a_first_address => 0,
	port_a_first_bit_number => 0,
	port_a_last_address => 511,
	port_a_logical_ram_depth => 258,
	port_a_logical_ram_width => 16,
	port_a_read_during_write_mode => "new_data_no_nbe_read",
	port_b_address_clear => "none",
	port_b_address_clock => "clock0",
	port_b_address_width => 9,
	port_b_data_out_clear => "none",
	port_b_data_out_clock => "none",
	port_b_data_width => 20,
	port_b_first_address => 0,
	port_b_first_bit_number => 0,
	port_b_last_address => 511,
	port_b_logical_ram_depth => 258,
	port_b_logical_ram_width => 16,
	port_b_read_during_write_mode => "new_data_no_nbe_read",
	port_b_read_enable_clock => "clock0",
	ram_block_type => "M20K")
-- pragma translate_on
PORT MAP (
	portawe => \TheI2sToPar|ValL~q\,
	portbre => VCC,
	clk0 => \iClk~inputCLKENA0_outclk\,
	portadatain => \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a4_PORTADATAIN_bus\,
	portaaddr => \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a4_PORTAADDR_bus\,
	portbaddr => \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a4_PORTBADDR_bus\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	portbdataout => \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a4_PORTBDATAOUT_bus\);

-- Location: MLABCELL_X15_Y61_N39
\TheRxFsk|Bandpasses:7:Bandpass0|Sample[-15]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-15]~0_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a0\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-15]~q\) # (\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\) ) 
-- ) # ( !\TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a0\ & ( (!\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-15]~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000101000001010010111110101111100001010000010100101111101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-15]~q\,
	datae => \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a0\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-15]~0_combout\);

-- Location: LABCELL_X18_Y63_N18
\TheRxFsk|Bandpasses:7:Bandpass0|Sample[-14]~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-14]~1_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a1\ ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & 
-- ( \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a1\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-14]~q\ ) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( 
-- !\TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a1\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-14]~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111000000000000000000001111000011111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-14]~q\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a1\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-14]~1_combout\);

-- Location: LABCELL_X19_Y63_N24
\TheRxFsk|Bandpasses:7:Bandpass0|Sample[-13]~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-13]~2_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a2\ ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & 
-- ( \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a2\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-13]~q\ ) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( 
-- !\TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a2\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-13]~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001100110011000000000000000000110011001100111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-13]~q\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a2\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-13]~2_combout\);

-- Location: LABCELL_X17_Y63_N0
\TheRxFsk|Bandpasses:7:Bandpass0|Sample[-12]~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-12]~3_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a3\ ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & 
-- ( \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a3\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-12]~q\ ) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( 
-- !\TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a3\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-12]~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001100110011000000000000000000110011001100111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-12]~q\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a3\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-12]~3_combout\);

-- Location: LABCELL_X17_Y63_N54
\TheRxFsk|Bandpasses:7:Bandpass0|Sample[-11]~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-11]~4_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a4\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\) # (\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-11]~q\) ) 
-- ) # ( !\TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a4\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-11]~q\ & !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011000000110000001100000011000000111111001111110011111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-11]~q\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a4\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-11]~4_combout\);

-- Location: LABCELL_X17_Y63_N27
\TheRxFsk|Bandpasses:7:Bandpass0|Sample[-10]~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-10]~5_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-10]~q\ & ( (!\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\) # (\TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a5\) 
-- ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-10]~q\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a5\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001010101000000000101010110101010111111111010101011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	datad => \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a5\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-10]~q\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-10]~5_combout\);

-- Location: LABCELL_X19_Y63_N36
\TheRxFsk|Bandpasses:7:Bandpass0|Sample[-9]~6\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-9]~6_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a6\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-9]~q\) # (\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\) ) ) 
-- # ( !\TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a6\ & ( (!\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-9]~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000101000001010000010100000101001011111010111110101111101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-9]~q\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a6\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-9]~6_combout\);

-- Location: LABCELL_X18_Y63_N39
\TheRxFsk|Bandpasses:7:Bandpass0|Sample[-8]~7\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-8]~7_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a7\ ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & 
-- ( \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a7\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-8]~q\ ) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( 
-- !\TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a7\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-8]~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111000000000000000000001111000011111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-8]~q\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a7\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-8]~7_combout\);

-- Location: MLABCELL_X15_Y63_N15
\TheRxFsk|Bandpasses:7:Bandpass0|Sample[-7]~8\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-7]~8_combout\ = (!\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ((\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-7]~q\))) # (\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & 
-- (\TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a8\))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001110100011101000111010001110100011101000111010001110100011101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a8\,
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-7]~q\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-7]~8_combout\);

-- Location: MLABCELL_X15_Y63_N21
\TheRxFsk|Bandpasses:7:Bandpass0|Sample[-6]~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-6]~9_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-6]~q\ & ( (!\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\) # (\TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a9\) ) 
-- ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-6]~q\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a9\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100000101000001010000010110101111101011111010111110101111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a9\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-6]~q\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-6]~9_combout\);

-- Location: LABCELL_X18_Y63_N30
\TheRxFsk|Bandpasses:7:Bandpass0|Sample[-5]~10\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-5]~10_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a10\ ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ 
-- & ( \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a10\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-5]~q\ ) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( 
-- !\TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a10\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-5]~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111000000000000000000001111000011111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-5]~q\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a10\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-5]~10_combout\);

-- Location: LABCELL_X16_Y63_N6
\TheRxFsk|Bandpasses:7:Bandpass0|Sample[-4]~11\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-4]~11_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-4]~q\ & ( \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a11\ ) ) # ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-4]~q\ & ( \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a11\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ ) ) ) # ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-4]~q\ 
-- & ( !\TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a11\ & ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000001111000011111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-4]~q\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a11\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-4]~11_combout\);

-- Location: LABCELL_X19_Y63_N30
\TheRxFsk|Bandpasses:7:Bandpass0|Sample[-3]~12\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-3]~12_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a12\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-3]~q\) # (\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\) ) 
-- ) # ( !\TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a12\ & ( (!\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-3]~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000101000001010000010100000101001011111010111110101111101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-3]~q\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a12\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-3]~12_combout\);

-- Location: LABCELL_X19_Y63_N3
\TheRxFsk|Bandpasses:7:Bandpass0|Sample[-2]~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-2]~13_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a13\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-2]~q\) # (\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\) ) 
-- ) # ( !\TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a13\ & ( (!\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-2]~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000010101010000000001010101001010101111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-2]~q\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a13\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-2]~13_combout\);

-- Location: LABCELL_X17_Y63_N24
\TheRxFsk|Bandpasses:7:Bandpass0|Sample[-1]~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-1]~14_combout\ = (!\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & (\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-1]~q\)) # (\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & 
-- ((\TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a14\)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000101001011111000010100101111100001010010111110000101001011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-1]~q\,
	datad => \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a14\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|Sample[-1]~14_combout\);

-- Location: LABCELL_X19_Y63_N21
\TheRxFsk|Bandpasses:7:Bandpass0|Sample[0]~15\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Sample[0]~15_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a15\ ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & 
-- ( \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a15\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[0]~DUPLICATE_q\ ) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( 
-- !\TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ram_block1a15\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[0]~DUPLICATE_q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010101010101000000000000000001010101010101011111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[0]~DUPLICATE_q\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass0|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a15\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|Sample[0]~15_combout\);

-- Location: DSP_X20_Y63_N0
\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8\ : cyclonev_mac
-- pragma translate_off
GENERIC MAP (
	accumulate_clock => "none",
	ax_clock => "none",
	ax_width => 18,
	ay_scan_in_clock => "none",
	ay_scan_in_width => 19,
	ay_use_scan_in => "false",
	az_clock => "none",
	bx_clock => "none",
	by_clock => "none",
	by_use_scan_in => "false",
	bz_clock => "none",
	coef_a_0 => 0,
	coef_a_1 => 0,
	coef_a_2 => 0,
	coef_a_3 => 0,
	coef_a_4 => 0,
	coef_a_5 => 0,
	coef_a_6 => 0,
	coef_a_7 => 0,
	coef_b_0 => 0,
	coef_b_1 => 0,
	coef_b_2 => 0,
	coef_b_3 => 0,
	coef_b_4 => 0,
	coef_b_5 => 0,
	coef_b_6 => 0,
	coef_b_7 => 0,
	coef_sel_a_clock => "none",
	coef_sel_b_clock => "none",
	delay_scan_out_ay => "false",
	delay_scan_out_by => "false",
	enable_double_accum => "false",
	load_const_clock => "none",
	load_const_value => 0,
	mode_sub_location => 0,
	negate_clock => "none",
	operand_source_max => "input",
	operand_source_may => "input",
	operand_source_mbx => "input",
	operand_source_mby => "input",
	operation_mode => "m18x18_full",
	output_clock => "none",
	preadder_subtract_a => "false",
	preadder_subtract_b => "false",
	result_a_width => 64,
	signed_max => "true",
	signed_may => "true",
	signed_mbx => "false",
	signed_mby => "false",
	sub_clock => "none",
	use_chainadder => "false")
-- pragma translate_on
PORT MAP (
	sub => GND,
	negate => GND,
	ax => \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_AX_bus\,
	ay => \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_AY_bus\,
	resulta => \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_RESULTA_bus\);

-- Location: LABCELL_X19_Y63_N54
\TheRxFsk|Bandpasses:7:Bandpass0|vAdd~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|vAdd~1_combout\ = ( !\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~14\ & ( !\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~9\ & ( (!\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~16\ & (!\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~18\ & 
-- (!\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~17\ & !\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~15\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1000000000000000000000000000000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~16\,
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~18\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~17\,
	datad => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~15\,
	datae => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~14\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~9\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|vAdd~1_combout\);

-- Location: LABCELL_X22_Y63_N6
\TheRxFsk|Bandpasses:7:Bandpass0|vAdd~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|vAdd~2_combout\ = ( !\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~10\ & ( !\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~11\ & ( (!\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~12\ & (!\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~8_resulta\ & 
-- !\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~21\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1000000010000000000000000000000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~12\,
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~8_resulta\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~21\,
	datae => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~10\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~11\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|vAdd~2_combout\);

-- Location: MLABCELL_X21_Y63_N54
\TheRxFsk|Bandpasses:7:Bandpass0|vAdd~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|vAdd~0_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass0|vAdd~2_combout\ & ( \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~19\ ) ) # ( !\TheRxFsk|Bandpasses:7:Bandpass0|vAdd~2_combout\ & ( \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~19\ ) 
-- ) # ( \TheRxFsk|Bandpasses:7:Bandpass0|vAdd~2_combout\ & ( !\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~19\ & ( (!\TheRxFsk|Bandpasses:7:Bandpass0|vAdd~1_combout\) # (((\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~13\) # (\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~22\)) 
-- # (\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~20\)) ) ) ) # ( !\TheRxFsk|Bandpasses:7:Bandpass0|vAdd~2_combout\ & ( !\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~19\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111111111111101111111111111111111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_vAdd~1_combout\,
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~20\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~22\,
	datad => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~13\,
	datae => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_vAdd~2_combout\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~19\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|vAdd~0_combout\);

-- Location: MLABCELL_X21_Y63_N0
\TheRxFsk|Bandpasses:7:Bandpass0|Add3~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add3~13_sumout\ = SUM(( (\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~39\ & \TheRxFsk|Bandpasses:7:Bandpass0|vAdd~0_combout\) ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~23\ ) + ( !VCC ))
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add3~14\ = CARRY(( (\TheRxFsk|Bandpasses:7:Bandpass0|Mult0~39\ & \TheRxFsk|Bandpasses:7:Bandpass0|vAdd~0_combout\) ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~23\ ) + ( !VCC ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000001010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~39\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~23\,
	datad => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_vAdd~0_combout\,
	cin => GND,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~13_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~14\);

-- Location: MLABCELL_X21_Y63_N3
\TheRxFsk|Bandpasses:7:Bandpass0|Add3~17\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add3~17_sumout\ = SUM(( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~24\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add3~14\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add3~18\ = CARRY(( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~24\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add3~14\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~24\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~14\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~17_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~18\);

-- Location: MLABCELL_X21_Y63_N6
\TheRxFsk|Bandpasses:7:Bandpass0|Add3~21\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add3~21_sumout\ = SUM(( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~25\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add3~18\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add3~22\ = CARRY(( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~25\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add3~18\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000110011001100110000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~25\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~18\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~21_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~22\);

-- Location: MLABCELL_X21_Y63_N9
\TheRxFsk|Bandpasses:7:Bandpass0|Add3~25\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add3~25_sumout\ = SUM(( \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~26\ ) + ( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add3~22\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add3~26\ = CARRY(( \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~26\ ) + ( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add3~22\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~26\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~22\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~25_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~26\);

-- Location: MLABCELL_X21_Y63_N12
\TheRxFsk|Bandpasses:7:Bandpass0|Add3~29\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add3~29_sumout\ = SUM(( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~27\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add3~26\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add3~30\ = CARRY(( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~27\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add3~26\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~27\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~26\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~29_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~30\);

-- Location: MLABCELL_X21_Y63_N15
\TheRxFsk|Bandpasses:7:Bandpass0|Add3~33\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add3~33_sumout\ = SUM(( \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~28\ ) + ( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add3~30\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add3~34\ = CARRY(( \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~28\ ) + ( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add3~30\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~28\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~30\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~33_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~34\);

-- Location: MLABCELL_X21_Y63_N18
\TheRxFsk|Bandpasses:7:Bandpass0|Add3~37\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add3~37_sumout\ = SUM(( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~29\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add3~34\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add3~38\ = CARRY(( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~29\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add3~34\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~29\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~34\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~37_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~38\);

-- Location: MLABCELL_X21_Y63_N21
\TheRxFsk|Bandpasses:7:Bandpass0|Add3~41\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add3~41_sumout\ = SUM(( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~30\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add3~38\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add3~42\ = CARRY(( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~30\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add3~38\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~30\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~38\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~41_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~42\);

-- Location: MLABCELL_X21_Y63_N24
\TheRxFsk|Bandpasses:7:Bandpass0|Add3~45\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add3~45_sumout\ = SUM(( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~31\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add3~42\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add3~46\ = CARRY(( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~31\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add3~42\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000110011001100110000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~31\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~42\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~45_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~46\);

-- Location: MLABCELL_X21_Y63_N27
\TheRxFsk|Bandpasses:7:Bandpass0|Add3~49\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add3~49_sumout\ = SUM(( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~32\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add3~46\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add3~50\ = CARRY(( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~32\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add3~46\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~32\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~46\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~49_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~50\);

-- Location: MLABCELL_X21_Y63_N30
\TheRxFsk|Bandpasses:7:Bandpass0|Add3~53\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add3~53_sumout\ = SUM(( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~33\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add3~50\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add3~54\ = CARRY(( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~33\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add3~50\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~33\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~50\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~53_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~54\);

-- Location: MLABCELL_X21_Y63_N33
\TheRxFsk|Bandpasses:7:Bandpass0|Add3~57\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add3~57_sumout\ = SUM(( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~34\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add3~54\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add3~58\ = CARRY(( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~34\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add3~54\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~34\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~54\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~57_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~58\);

-- Location: MLABCELL_X21_Y63_N36
\TheRxFsk|Bandpasses:7:Bandpass0|Add3~61\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add3~61_sumout\ = SUM(( \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~35\ ) + ( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add3~58\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add3~62\ = CARRY(( \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~35\ ) + ( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add3~58\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~35\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~58\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~61_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~62\);

-- Location: MLABCELL_X21_Y63_N39
\TheRxFsk|Bandpasses:7:Bandpass0|Add3~65\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add3~65_sumout\ = SUM(( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~36\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add3~62\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add3~66\ = CARRY(( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~36\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add3~62\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~36\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~62\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~65_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~66\);

-- Location: MLABCELL_X21_Y63_N42
\TheRxFsk|Bandpasses:7:Bandpass0|Add3~69\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add3~69_sumout\ = SUM(( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~37\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add3~66\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add3~70\ = CARRY(( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~37\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add3~66\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~37\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~66\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~69_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~70\);

-- Location: MLABCELL_X21_Y63_N45
\TheRxFsk|Bandpasses:7:Bandpass0|Add3~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add3~9_sumout\ = SUM(( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~38\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add3~70\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add3~10\ = CARRY(( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~38\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add3~70\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~38\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~70\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~9_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~10\);

-- Location: MLABCELL_X21_Y63_N48
\TheRxFsk|Bandpasses:7:Bandpass0|Add3~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add3~5_sumout\ = SUM(( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~39\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add3~10\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add3~6\ = CARRY(( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~39\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add3~10\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~39\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~10\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~5_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~6\);

-- Location: MLABCELL_X21_Y63_N51
\TheRxFsk|Bandpasses:7:Bandpass0|Add3~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add3~1_sumout\ = SUM(( VCC ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Mult0~39\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add3~6\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000101010101010101000000000000000001111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Mult0~39\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~6\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~1_sumout\);

-- Location: MLABCELL_X21_Y64_N0
\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[0]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[0]~0_combout\ = ( !\TheRxFsk|Bandpasses:7:Bandpass0|Add3~1_sumout\ )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111111111111111111111111111100000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add3~1_sumout\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[0]~0_combout\);

-- Location: FF_X21_Y64_N1
\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[0]~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed\(0));

-- Location: FF_X21_Y63_N46
\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_NEW_REG68\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~9_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM69\);

-- Location: FF_X21_Y63_N43
\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-1]_NEW_REG96\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~69_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-1]_OTERM97\);

-- Location: FF_X21_Y63_N49
\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_NEW_REG66\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~5_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM67\);

-- Location: FF_X21_Y63_N53
\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_NEW_REG64\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~1_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM65\);

-- Location: LABCELL_X22_Y63_N15
\TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-1]~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-1]~14_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM65\ & ( ((\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM67\) # 
-- (\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-1]_OTERM97\)) # (\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM69\) ) ) # ( !\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM65\ & ( 
-- (\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM69\ & (\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-1]_OTERM97\ & \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM67\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000100000001011111110111111100000001000000010111111101111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM69\,
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-1]_OTERM97\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM67\,
	datae => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM65\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-1]~14_combout\);

-- Location: FF_X21_Y63_N40
\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-2]_NEW_REG102\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~65_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-2]_OTERM103\);

-- Location: LABCELL_X22_Y63_N21
\TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-2]~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-2]~13_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-2]_OTERM103\ & ( ((\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM69\ & 
-- \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM67\)) # (\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM65\) ) ) # ( !\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-2]_OTERM103\ & ( 
-- (\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM65\ & ((\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM67\) # (\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM69\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000011100000111000001110000011100011111000111110001111100011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM69\,
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM67\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM65\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-2]_OTERM103\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-2]~13_combout\);

-- Location: LABCELL_X19_Y64_N45
\TheRxFsk|Bandpasses:7:Bandpass0|Add4~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add4~5_sumout\ = SUM(( \TheRxFsk|Bandpasses:7:Bandpass0|Sum\(0) ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed\(0) ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add4~66\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add4~6\ = CARRY(( \TheRxFsk|Bandpasses:7:Bandpass0|Sum\(0) ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed\(0) ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add4~66\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111110000000000000000000000000101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum\(0),
	dataf => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed\(0),
	cin => \TheRxFsk|Bandpasses:7:Bandpass0|Add4~66\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass0|Add4~5_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass0|Add4~6\);

-- Location: FF_X21_Y63_N37
\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-3]_NEW_REG108\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~61_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-3]_OTERM109\);

-- Location: LABCELL_X22_Y63_N18
\TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-3]~12\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-3]~12_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-3]_OTERM109\ & ( ((\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM69\ & 
-- \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM67\)) # (\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM65\) ) ) # ( !\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-3]_OTERM109\ & ( 
-- (\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM65\ & ((\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM67\) # (\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM69\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001110111000000000111011100010001111111110001000111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM69\,
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM67\,
	datad => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM65\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-3]_OTERM109\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-3]~12_combout\);

-- Location: FF_X21_Y63_N34
\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-4]_NEW_REG114\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~57_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-4]_OTERM115\);

-- Location: LABCELL_X22_Y63_N51
\TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-4]~11\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-4]~11_combout\ = (!\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM69\ & (\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM65\ & 
-- ((\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-4]_OTERM115\) # (\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM67\)))) # (\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM69\ & 
-- (((\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM67\ & \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-4]_OTERM115\)) # (\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM65\)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000101111111000000010111111100000001011111110000000101111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM69\,
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM67\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-4]_OTERM115\,
	datad => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM65\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-4]~11_combout\);

-- Location: FF_X21_Y63_N31
\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-5]_NEW_REG120\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~53_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-5]_OTERM121\);

-- Location: LABCELL_X22_Y63_N48
\TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-5]~10\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-5]~10_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-5]_OTERM121\ & ( ((\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM69\ & 
-- \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM67\)) # (\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM65\) ) ) # ( !\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-5]_OTERM121\ & ( 
-- (\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM65\ & ((\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM67\) # (\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM69\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001110111000000000111011100010001111111110001000111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM69\,
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM67\,
	datad => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM65\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-5]_OTERM121\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-5]~10_combout\);

-- Location: FF_X21_Y63_N28
\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-6]_NEW_REG126\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~49_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-6]_OTERM127\);

-- Location: LABCELL_X22_Y63_N33
\TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-6]~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-6]~9_combout\ = (!\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM69\ & (\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM65\ & 
-- ((\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-6]_OTERM127\) # (\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM67\)))) # (\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM69\ & 
-- (((\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM67\ & \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-6]_OTERM127\)) # (\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM65\)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000011100011111000001110001111100000111000111110000011100011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM69\,
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM67\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM65\,
	datad => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-6]_OTERM127\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-6]~9_combout\);

-- Location: FF_X21_Y63_N25
\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-7]_NEW_REG132\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~45_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-7]_OTERM133\);

-- Location: LABCELL_X22_Y63_N30
\TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-7]~8\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-7]~8_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-7]_OTERM133\ & ( ((\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM69\ & 
-- \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM67\)) # (\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM65\) ) ) # ( !\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-7]_OTERM133\ & ( 
-- (\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM65\ & ((\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM67\) # (\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM69\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001110111000000000111011100010001111111110001000111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM69\,
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM67\,
	datad => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM65\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-7]_OTERM133\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-7]~8_combout\);

-- Location: FF_X21_Y63_N22
\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-8]_NEW_REG138\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~41_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-8]_OTERM139\);

-- Location: LABCELL_X22_Y63_N39
\TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-8]~7\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-8]~7_combout\ = (!\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM69\ & (\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM65\ & 
-- ((\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-8]_OTERM139\) # (\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM67\)))) # (\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM69\ & 
-- (((\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM67\ & \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-8]_OTERM139\)) # (\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM65\)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000011100011111000001110001111100000111000111110000011100011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM69\,
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM67\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM65\,
	datad => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-8]_OTERM139\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-8]~7_combout\);

-- Location: FF_X21_Y63_N19
\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-9]_NEW_REG144\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~37_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-9]_OTERM145\);

-- Location: LABCELL_X22_Y63_N36
\TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-9]~6\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-9]~6_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-9]_OTERM145\ & ( ((\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM69\ & 
-- \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM67\)) # (\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM65\) ) ) # ( !\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-9]_OTERM145\ & ( 
-- (\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM65\ & ((\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM67\) # (\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM69\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001110111000000000111011100010001111111110001000111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM69\,
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM67\,
	datad => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM65\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-9]_OTERM145\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-9]~6_combout\);

-- Location: FF_X21_Y63_N16
\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-10]_NEW_REG150\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~33_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-10]_OTERM151\);

-- Location: LABCELL_X22_Y63_N45
\TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-10]~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-10]~5_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-10]_OTERM151\ & ( ((\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM69\ & 
-- \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM67\)) # (\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM65\) ) ) # ( !\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-10]_OTERM151\ & ( 
-- (\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM65\ & ((\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM67\) # (\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM69\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000011100000111000001110000011100011111000111110001111100011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM69\,
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM67\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM65\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-10]_OTERM151\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-10]~5_combout\);

-- Location: FF_X21_Y63_N13
\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-11]_NEW_REG156\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~29_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-11]_OTERM157\);

-- Location: LABCELL_X22_Y63_N42
\TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-11]~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-11]~4_combout\ = (!\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM69\ & (\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM65\ & 
-- ((\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-11]_OTERM157\) # (\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM67\)))) # (\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM69\ & 
-- (((\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM67\ & \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-11]_OTERM157\)) # (\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM65\)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000101111111000000010111111100000001011111110000000101111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM69\,
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM67\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-11]_OTERM157\,
	datad => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM65\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-11]~4_combout\);

-- Location: FF_X21_Y63_N10
\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-12]_NEW_REG162\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~25_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-12]_OTERM163\);

-- Location: LABCELL_X22_Y63_N3
\TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-12]~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-12]~3_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-12]_OTERM163\ & ( ((\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM69\ & 
-- \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM67\)) # (\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM65\) ) ) # ( !\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-12]_OTERM163\ & ( 
-- (\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM65\ & ((\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM67\) # (\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM69\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001001100010011001101110011011100010011000100110011011100110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM69\,
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM65\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM67\,
	datae => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-12]_OTERM163\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-12]~3_combout\);

-- Location: FF_X21_Y63_N7
\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-13]_NEW_REG168\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~21_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-13]_OTERM169\);

-- Location: LABCELL_X22_Y63_N54
\TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-13]~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-13]~2_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM65\ & ( \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM69\ ) ) # ( 
-- !\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM65\ & ( \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM69\ & ( (\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM67\ & 
-- \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-13]_OTERM169\) ) ) ) # ( \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM65\ & ( !\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM69\ & ( 
-- (\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-13]_OTERM169\) # (\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM67\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000001111110011111100000011000000111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM67\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-13]_OTERM169\,
	datae => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM65\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM69\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-13]~2_combout\);

-- Location: FF_X21_Y63_N4
\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-14]_NEW_REG174\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~17_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-14]_OTERM175\);

-- Location: LABCELL_X23_Y63_N27
\TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-14]~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-14]~1_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM65\ & ( \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-14]_OTERM175\ ) ) # ( 
-- !\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM65\ & ( \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-14]_OTERM175\ & ( (\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM69\ & 
-- \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM67\) ) ) ) # ( \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM65\ & ( !\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-14]_OTERM175\ & ( 
-- (\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM67\) # (\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM69\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000001111110011111100000011000000111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM69\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM67\,
	datae => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM65\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-14]_OTERM175\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-14]~1_combout\);

-- Location: FF_X21_Y63_N1
\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_NEW_REG70\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass0|Add3~13_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM71\);

-- Location: LABCELL_X22_Y63_N27
\TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-15]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-15]~0_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM65\ & ( \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM69\ ) ) # ( 
-- !\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM65\ & ( \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM69\ & ( (\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM71\ & 
-- \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM67\) ) ) ) # ( \TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM65\ & ( !\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM69\ & ( 
-- (\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM67\) # (\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed[-15]_OTERM71\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000001111110011111100000011000000111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM71\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM67\,
	datae => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM65\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed[-15]_OTERM69\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-15]~0_combout\);

-- Location: LABCELL_X18_Y64_N42
\TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-15]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-15]~0_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-15]~0_combout\ & ( (!\TheRxFsk|Bandpasses:7:Bandpass0|Add4~5_sumout\ & (\TheRxFsk|Bandpasses:7:Bandpass0|Add4~1_sumout\ & 
-- !\TheRxFsk|Bandpasses:7:Bandpass0|Sum[-15]~q\)) # (\TheRxFsk|Bandpasses:7:Bandpass0|Add4~5_sumout\ & ((!\TheRxFsk|Bandpasses:7:Bandpass0|Sum[-15]~q\) # (\TheRxFsk|Bandpasses:7:Bandpass0|Add4~1_sumout\))) ) ) # ( 
-- !\TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-15]~0_combout\ & ( (!\TheRxFsk|Bandpasses:7:Bandpass0|Add4~5_sumout\ & (\TheRxFsk|Bandpasses:7:Bandpass0|Add4~1_sumout\ & \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-15]~q\)) # 
-- (\TheRxFsk|Bandpasses:7:Bandpass0|Add4~5_sumout\ & ((\TheRxFsk|Bandpasses:7:Bandpass0|Sum[-15]~q\) # (\TheRxFsk|Bandpasses:7:Bandpass0|Add4~1_sumout\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000101110111000100010111011101110111000100010111011100010001",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~5_sumout\,
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~1_sumout\,
	datad => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-15]~q\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResult[-15]~0_combout\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-15]~0_combout\);

-- Location: FF_X21_Y64_N23
\TheRxFsk|Bandpasses:7:Bandpass0|R.SumState.SumValid\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	asdata => \TheRxFsk|Bandpasses:7:Bandpass0|R.SumState.SumWait2~q\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass0|R.SumState.SumValid~q\);

-- Location: MLABCELL_X21_Y64_N33
\TheRxFsk|Bandpasses:7:Bandpass0|Selector0~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Selector0~0_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass0|R.SumState.Idle~q\ & ( \TheI2sToPar|ValL~q\ & ( !\TheRxFsk|Bandpasses:7:Bandpass0|R.SumState.SumValid~q\ ) ) ) # ( 
-- !\TheRxFsk|Bandpasses:7:Bandpass0|R.SumState.Idle~q\ & ( \TheI2sToPar|ValL~q\ & ( !\TheRxFsk|Bandpasses:7:Bandpass0|R.SumState.SumValid~q\ ) ) ) # ( \TheRxFsk|Bandpasses:7:Bandpass0|R.SumState.Idle~q\ & ( !\TheI2sToPar|ValL~q\ & ( 
-- !\TheRxFsk|Bandpasses:7:Bandpass0|R.SumState.SumValid~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111110000000011111111000000001111111100000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_R.SumState.SumValid~q\,
	datae => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_R.SumState.Idle~q\,
	dataf => \TheI2sToPar|ALT_INV_ValL~q\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|Selector0~0_combout\);

-- Location: FF_X21_Y64_N35
\TheRxFsk|Bandpasses:7:Bandpass0|R.SumState.Idle\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass0|Selector0~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass0|R.SumState.Idle~q\);

-- Location: MLABCELL_X21_Y64_N48
\TheRxFsk|Bandpasses:7:Bandpass0|Selector1~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Selector1~0_combout\ = ( \TheI2sToPar|ValL~q\ & ( !\TheRxFsk|Bandpasses:7:Bandpass0|R.SumState.Idle~q\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000010101010101010101010101010101010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_R.SumState.Idle~q\,
	dataf => \TheI2sToPar|ALT_INV_ValL~q\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|Selector1~0_combout\);

-- Location: FF_X21_Y64_N49
\TheRxFsk|Bandpasses:7:Bandpass0|R.SumState.SumEnable\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass0|Selector1~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass0|R.SumState.SumEnable~q\);

-- Location: MLABCELL_X21_Y64_N12
\TheRxFsk|Bandpasses:7:Bandpass0|Selector2~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Selector2~0_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass0|R.SumState.SumEnable~q\ ) # ( !\TheRxFsk|Bandpasses:7:Bandpass0|R.SumState.SumEnable~q\ & ( (\TheRxFsk|Bandpasses:7:Bandpass0|R.SumState.SumSelect~q\ & 
-- ((!\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~0_combout\) # (!\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~1_combout\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011101110000000001110111011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:11:Bandpass1|ALT_INV_Equal1~0_combout\,
	datab => \TheRxFsk|Bandpasses:11:Bandpass1|ALT_INV_Equal1~1_combout\,
	datad => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_R.SumState.SumSelect~q\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_R.SumState.SumEnable~q\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|Selector2~0_combout\);

-- Location: FF_X21_Y64_N13
\TheRxFsk|Bandpasses:7:Bandpass0|R.SumState.SumSelect\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass0|Selector2~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass0|R.SumState.SumSelect~q\);

-- Location: MLABCELL_X21_Y64_N15
\TheRxFsk|Bandpasses:7:Bandpass0|Selector3~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Selector3~0_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass0|R.SumState.SumSelect~q\ & ( (\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~0_combout\ & \TheRxFsk|Bandpasses:11:Bandpass1|Equal1~1_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000010001000100010001000100010001",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:11:Bandpass1|ALT_INV_Equal1~0_combout\,
	datab => \TheRxFsk|Bandpasses:11:Bandpass1|ALT_INV_Equal1~1_combout\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_R.SumState.SumSelect~q\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|Selector3~0_combout\);

-- Location: FF_X21_Y64_N17
\TheRxFsk|Bandpasses:7:Bandpass0|R.SumState.SumWait1\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass0|Selector3~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass0|R.SumState.SumWait1~q\);

-- Location: FF_X21_Y64_N47
\TheRxFsk|Bandpasses:7:Bandpass0|R.SumState.SumWait2\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	asdata => \TheRxFsk|Bandpasses:7:Bandpass0|R.SumState.SumWait1~q\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass0|R.SumState.SumWait2~q\);

-- Location: MLABCELL_X21_Y64_N57
\TheRxFsk|Bandpasses:7:Bandpass0|Selector6~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Selector6~0_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass0|R.SelSumUp~q\ & ( \TheRxFsk|Bandpasses:7:Bandpass0|R.SumState.SumEnable~q\ ) ) # ( !\TheRxFsk|Bandpasses:7:Bandpass0|R.SelSumUp~q\ & ( 
-- \TheRxFsk|Bandpasses:7:Bandpass0|R.SumState.SumEnable~q\ ) ) # ( \TheRxFsk|Bandpasses:7:Bandpass0|R.SelSumUp~q\ & ( !\TheRxFsk|Bandpasses:7:Bandpass0|R.SumState.SumEnable~q\ & ( !\TheRxFsk|Bandpasses:7:Bandpass0|R.SumState.SumWait2~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000110011001100110011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_R.SumState.SumWait2~q\,
	datae => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_R.SelSumUp~q\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_R.SumState.SumEnable~q\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|Selector6~0_combout\);

-- Location: FF_X21_Y64_N59
\TheRxFsk|Bandpasses:7:Bandpass0|R.SelSumUp\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass0|Selector6~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass0|R.SelSumUp~q\);

-- Location: FF_X21_Y64_N34
\TheRxFsk|Bandpasses:7:Bandpass0|R.SumState.Idle~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass0|Selector0~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass0|R.SumState.Idle~DUPLICATE_q\);

-- Location: LABCELL_X18_Y64_N21
\TheRxFsk|Bandpasses:7:Bandpass0|Selector7~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Selector7~0_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass0|R.EnableSumUp~q\ & ( \TheI2sToPar|ValL~q\ & ( (!\TheRxFsk|Bandpasses:7:Bandpass0|R.SumState.Idle~DUPLICATE_q\) # 
-- (!\TheRxFsk|Bandpasses:7:Bandpass0|R.SumState.SumWait2~q\) ) ) ) # ( !\TheRxFsk|Bandpasses:7:Bandpass0|R.EnableSumUp~q\ & ( \TheI2sToPar|ValL~q\ & ( !\TheRxFsk|Bandpasses:7:Bandpass0|R.SumState.Idle~DUPLICATE_q\ ) ) ) # ( 
-- \TheRxFsk|Bandpasses:7:Bandpass0|R.EnableSumUp~q\ & ( !\TheI2sToPar|ValL~q\ & ( (!\TheRxFsk|Bandpasses:7:Bandpass0|R.SumState.Idle~DUPLICATE_q\) # (!\TheRxFsk|Bandpasses:7:Bandpass0|R.SumState.SumWait2~q\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111110101111101010101010101010101111101011111010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_R.SumState.Idle~DUPLICATE_q\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_R.SumState.SumWait2~q\,
	datae => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_R.EnableSumUp~q\,
	dataf => \TheI2sToPar|ALT_INV_ValL~q\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|Selector7~0_combout\);

-- Location: FF_X18_Y64_N23
\TheRxFsk|Bandpasses:7:Bandpass0|R.EnableSumUp\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass0|Selector7~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass0|R.EnableSumUp~q\);

-- Location: FF_X18_Y64_N43
\TheRxFsk|Bandpasses:7:Bandpass0|Sum[-15]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-15]~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:7:Bandpass0|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-15]~q\);

-- Location: LABCELL_X19_Y64_N0
\TheRxFsk|Bandpasses:7:Bandpass0|Add4~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add4~10\ = CARRY(( \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-15]~q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-15]~0_combout\ ) + ( !VCC ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111110000000000000000000000000011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-15]~q\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResult[-15]~0_combout\,
	cin => GND,
	cout => \TheRxFsk|Bandpasses:7:Bandpass0|Add4~10\);

-- Location: LABCELL_X19_Y64_N3
\TheRxFsk|Bandpasses:7:Bandpass0|Add4~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add4~13_sumout\ = SUM(( \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-14]~q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-14]~1_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add4~10\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add4~14\ = CARRY(( \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-14]~q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-14]~1_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add4~10\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000101010101010101000000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResult[-14]~1_combout\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-14]~q\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass0|Add4~10\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass0|Add4~13_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass0|Add4~14\);

-- Location: LABCELL_X19_Y64_N54
\TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-14]~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-14]~1_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass0|Add4~1_sumout\ & ( (\TheRxFsk|Bandpasses:7:Bandpass0|Add4~13_sumout\) # (\TheRxFsk|Bandpasses:7:Bandpass0|Add4~5_sumout\) ) ) # ( 
-- !\TheRxFsk|Bandpasses:7:Bandpass0|Add4~1_sumout\ & ( (\TheRxFsk|Bandpasses:7:Bandpass0|Add4~5_sumout\ & \TheRxFsk|Bandpasses:7:Bandpass0|Add4~13_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100000011000000110000001100111111001111110011111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~5_sumout\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~13_sumout\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~1_sumout\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-14]~1_combout\);

-- Location: FF_X19_Y64_N55
\TheRxFsk|Bandpasses:7:Bandpass0|Sum[-14]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-14]~1_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:7:Bandpass0|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-14]~q\);

-- Location: LABCELL_X19_Y64_N6
\TheRxFsk|Bandpasses:7:Bandpass0|Add4~17\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add4~17_sumout\ = SUM(( \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-13]~q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-13]~2_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add4~14\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add4~18\ = CARRY(( \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-13]~q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-13]~2_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add4~14\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-13]~q\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResult[-13]~2_combout\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass0|Add4~14\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass0|Add4~17_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass0|Add4~18\);

-- Location: LABCELL_X18_Y64_N48
\TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-13]~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-13]~2_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass0|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:7:Bandpass0|Add4~17_sumout\) # (\TheRxFsk|Bandpasses:7:Bandpass0|Add4~1_sumout\) ) ) # ( 
-- !\TheRxFsk|Bandpasses:7:Bandpass0|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:7:Bandpass0|Add4~1_sumout\ & \TheRxFsk|Bandpasses:7:Bandpass0|Add4~17_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100000011000000110000001100111111001111110011111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~1_sumout\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~17_sumout\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~5_sumout\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-13]~2_combout\);

-- Location: FF_X18_Y64_N49
\TheRxFsk|Bandpasses:7:Bandpass0|Sum[-13]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-13]~2_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:7:Bandpass0|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-13]~q\);

-- Location: LABCELL_X19_Y64_N9
\TheRxFsk|Bandpasses:7:Bandpass0|Add4~21\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add4~21_sumout\ = SUM(( \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-12]~3_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-12]~q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add4~18\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add4~22\ = CARRY(( \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-12]~3_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-12]~q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add4~18\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111110000000000000000000000000101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResult[-12]~3_combout\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-12]~q\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass0|Add4~18\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass0|Add4~21_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass0|Add4~22\);

-- Location: LABCELL_X18_Y64_N51
\TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-12]~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-12]~3_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass0|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:7:Bandpass0|Add4~21_sumout\) # (\TheRxFsk|Bandpasses:7:Bandpass0|Add4~1_sumout\) ) ) # ( 
-- !\TheRxFsk|Bandpasses:7:Bandpass0|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:7:Bandpass0|Add4~1_sumout\ & \TheRxFsk|Bandpasses:7:Bandpass0|Add4~21_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000110011000000000011001100110011111111110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~1_sumout\,
	datad => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~21_sumout\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~5_sumout\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-12]~3_combout\);

-- Location: FF_X18_Y64_N52
\TheRxFsk|Bandpasses:7:Bandpass0|Sum[-12]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-12]~3_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:7:Bandpass0|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-12]~q\);

-- Location: LABCELL_X19_Y64_N12
\TheRxFsk|Bandpasses:7:Bandpass0|Add4~25\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add4~25_sumout\ = SUM(( \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-11]~q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-11]~4_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add4~22\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add4~26\ = CARRY(( \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-11]~q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-11]~4_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add4~22\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResult[-11]~4_combout\,
	datad => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-11]~q\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass0|Add4~22\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass0|Add4~25_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass0|Add4~26\);

-- Location: LABCELL_X18_Y64_N54
\TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-11]~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-11]~4_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass0|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:7:Bandpass0|Add4~25_sumout\) # (\TheRxFsk|Bandpasses:7:Bandpass0|Add4~1_sumout\) ) ) # ( 
-- !\TheRxFsk|Bandpasses:7:Bandpass0|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:7:Bandpass0|Add4~1_sumout\ & \TheRxFsk|Bandpasses:7:Bandpass0|Add4~25_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100000011000000110000001100111111001111110011111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~1_sumout\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~25_sumout\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~5_sumout\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-11]~4_combout\);

-- Location: FF_X18_Y64_N55
\TheRxFsk|Bandpasses:7:Bandpass0|Sum[-11]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-11]~4_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:7:Bandpass0|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-11]~q\);

-- Location: LABCELL_X19_Y64_N15
\TheRxFsk|Bandpasses:7:Bandpass0|Add4~29\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add4~29_sumout\ = SUM(( \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-10]~q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-10]~5_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add4~26\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add4~30\ = CARRY(( \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-10]~q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-10]~5_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add4~26\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000101010101010101000000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResult[-10]~5_combout\,
	datad => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-10]~q\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass0|Add4~26\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass0|Add4~29_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass0|Add4~30\);

-- Location: LABCELL_X18_Y64_N57
\TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-10]~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-10]~5_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass0|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:7:Bandpass0|Add4~29_sumout\) # (\TheRxFsk|Bandpasses:7:Bandpass0|Add4~1_sumout\) ) ) # ( 
-- !\TheRxFsk|Bandpasses:7:Bandpass0|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:7:Bandpass0|Add4~1_sumout\ & \TheRxFsk|Bandpasses:7:Bandpass0|Add4~29_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000110011000000000011001100110011111111110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~1_sumout\,
	datad => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~29_sumout\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~5_sumout\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-10]~5_combout\);

-- Location: FF_X18_Y64_N58
\TheRxFsk|Bandpasses:7:Bandpass0|Sum[-10]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-10]~5_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:7:Bandpass0|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-10]~q\);

-- Location: LABCELL_X19_Y64_N18
\TheRxFsk|Bandpasses:7:Bandpass0|Add4~33\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add4~33_sumout\ = SUM(( \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-9]~6_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-9]~q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add4~30\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add4~34\ = CARRY(( \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-9]~6_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-9]~q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add4~30\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000110011001100110000000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-9]~q\,
	datad => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResult[-9]~6_combout\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass0|Add4~30\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass0|Add4~33_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass0|Add4~34\);

-- Location: LABCELL_X18_Y64_N0
\TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-9]~6\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-9]~6_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass0|Add4~33_sumout\ & ( (\TheRxFsk|Bandpasses:7:Bandpass0|Add4~1_sumout\) # (\TheRxFsk|Bandpasses:7:Bandpass0|Add4~5_sumout\) ) ) # ( 
-- !\TheRxFsk|Bandpasses:7:Bandpass0|Add4~33_sumout\ & ( (\TheRxFsk|Bandpasses:7:Bandpass0|Add4~5_sumout\ & \TheRxFsk|Bandpasses:7:Bandpass0|Add4~1_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000100010001000100010001000101110111011101110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~5_sumout\,
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~1_sumout\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~33_sumout\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-9]~6_combout\);

-- Location: FF_X18_Y64_N1
\TheRxFsk|Bandpasses:7:Bandpass0|Sum[-9]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-9]~6_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:7:Bandpass0|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-9]~q\);

-- Location: LABCELL_X19_Y64_N21
\TheRxFsk|Bandpasses:7:Bandpass0|Add4~37\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add4~37_sumout\ = SUM(( \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-8]~q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-8]~7_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add4~34\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add4~38\ = CARRY(( \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-8]~q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-8]~7_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add4~34\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111110000000000000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-8]~q\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResult[-8]~7_combout\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass0|Add4~34\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass0|Add4~37_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass0|Add4~38\);

-- Location: LABCELL_X18_Y64_N3
\TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-8]~7\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-8]~7_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass0|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:7:Bandpass0|Add4~37_sumout\) # (\TheRxFsk|Bandpasses:7:Bandpass0|Add4~1_sumout\) ) ) # ( 
-- !\TheRxFsk|Bandpasses:7:Bandpass0|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:7:Bandpass0|Add4~1_sumout\ & \TheRxFsk|Bandpasses:7:Bandpass0|Add4~37_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000110011000000000011001100110011111111110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~1_sumout\,
	datad => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~37_sumout\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~5_sumout\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-8]~7_combout\);

-- Location: FF_X18_Y64_N4
\TheRxFsk|Bandpasses:7:Bandpass0|Sum[-8]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-8]~7_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:7:Bandpass0|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-8]~q\);

-- Location: LABCELL_X19_Y64_N24
\TheRxFsk|Bandpasses:7:Bandpass0|Add4~41\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add4~41_sumout\ = SUM(( \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-7]~DUPLICATE_q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-7]~8_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add4~38\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add4~42\ = CARRY(( \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-7]~DUPLICATE_q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-7]~8_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add4~38\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111110000000000000000000000000101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-7]~DUPLICATE_q\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResult[-7]~8_combout\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass0|Add4~38\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass0|Add4~41_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass0|Add4~42\);

-- Location: LABCELL_X18_Y64_N6
\TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-7]~8\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-7]~8_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass0|Add4~41_sumout\ & ( (\TheRxFsk|Bandpasses:7:Bandpass0|Add4~1_sumout\) # (\TheRxFsk|Bandpasses:7:Bandpass0|Add4~5_sumout\) ) ) # ( 
-- !\TheRxFsk|Bandpasses:7:Bandpass0|Add4~41_sumout\ & ( (\TheRxFsk|Bandpasses:7:Bandpass0|Add4~5_sumout\ & \TheRxFsk|Bandpasses:7:Bandpass0|Add4~1_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000100010001000100010001000101110111011101110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~5_sumout\,
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~1_sumout\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~41_sumout\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-7]~8_combout\);

-- Location: FF_X18_Y64_N7
\TheRxFsk|Bandpasses:7:Bandpass0|Sum[-7]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-7]~8_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:7:Bandpass0|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-7]~DUPLICATE_q\);

-- Location: LABCELL_X19_Y64_N27
\TheRxFsk|Bandpasses:7:Bandpass0|Add4~45\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add4~45_sumout\ = SUM(( \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-6]~q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-6]~9_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add4~42\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add4~46\ = CARRY(( \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-6]~q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-6]~9_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add4~42\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000110011001100110000000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResult[-6]~9_combout\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-6]~q\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass0|Add4~42\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass0|Add4~45_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass0|Add4~46\);

-- Location: LABCELL_X18_Y64_N9
\TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-6]~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-6]~9_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass0|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:7:Bandpass0|Add4~45_sumout\) # (\TheRxFsk|Bandpasses:7:Bandpass0|Add4~1_sumout\) ) ) # ( 
-- !\TheRxFsk|Bandpasses:7:Bandpass0|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:7:Bandpass0|Add4~1_sumout\ & \TheRxFsk|Bandpasses:7:Bandpass0|Add4~45_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000110011000000000011001100110011111111110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~1_sumout\,
	datad => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~45_sumout\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~5_sumout\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-6]~9_combout\);

-- Location: FF_X18_Y64_N10
\TheRxFsk|Bandpasses:7:Bandpass0|Sum[-6]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-6]~9_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:7:Bandpass0|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-6]~q\);

-- Location: LABCELL_X19_Y64_N30
\TheRxFsk|Bandpasses:7:Bandpass0|Add4~49\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add4~49_sumout\ = SUM(( \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-5]~q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-5]~10_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add4~46\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add4~50\ = CARRY(( \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-5]~q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-5]~10_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add4~46\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111110000000000000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-5]~q\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResult[-5]~10_combout\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass0|Add4~46\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass0|Add4~49_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass0|Add4~50\);

-- Location: LABCELL_X18_Y64_N12
\TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-5]~10\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-5]~10_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass0|Add4~49_sumout\ & ( (\TheRxFsk|Bandpasses:7:Bandpass0|Add4~1_sumout\) # (\TheRxFsk|Bandpasses:7:Bandpass0|Add4~5_sumout\) ) ) # ( 
-- !\TheRxFsk|Bandpasses:7:Bandpass0|Add4~49_sumout\ & ( (\TheRxFsk|Bandpasses:7:Bandpass0|Add4~5_sumout\ & \TheRxFsk|Bandpasses:7:Bandpass0|Add4~1_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000100010001000100010001000101110111011101110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~5_sumout\,
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~1_sumout\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~49_sumout\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-5]~10_combout\);

-- Location: FF_X18_Y64_N13
\TheRxFsk|Bandpasses:7:Bandpass0|Sum[-5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-5]~10_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:7:Bandpass0|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-5]~q\);

-- Location: LABCELL_X19_Y64_N33
\TheRxFsk|Bandpasses:7:Bandpass0|Add4~53\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add4~53_sumout\ = SUM(( \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-4]~q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-4]~11_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add4~50\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add4~54\ = CARRY(( \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-4]~q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-4]~11_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add4~50\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000101010101010101000000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResult[-4]~11_combout\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-4]~q\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass0|Add4~50\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass0|Add4~53_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass0|Add4~54\);

-- Location: LABCELL_X18_Y64_N15
\TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-4]~11\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-4]~11_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass0|Add4~53_sumout\ & ( (\TheRxFsk|Bandpasses:7:Bandpass0|Add4~1_sumout\) # (\TheRxFsk|Bandpasses:7:Bandpass0|Add4~5_sumout\) ) ) # ( 
-- !\TheRxFsk|Bandpasses:7:Bandpass0|Add4~53_sumout\ & ( (\TheRxFsk|Bandpasses:7:Bandpass0|Add4~5_sumout\ & \TheRxFsk|Bandpasses:7:Bandpass0|Add4~1_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000100010001000100010001000101110111011101110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~5_sumout\,
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~1_sumout\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~53_sumout\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-4]~11_combout\);

-- Location: FF_X18_Y64_N16
\TheRxFsk|Bandpasses:7:Bandpass0|Sum[-4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-4]~11_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:7:Bandpass0|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-4]~q\);

-- Location: LABCELL_X19_Y64_N36
\TheRxFsk|Bandpasses:7:Bandpass0|Add4~57\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add4~57_sumout\ = SUM(( \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-3]~12_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-3]~q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add4~54\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add4~58\ = CARRY(( \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-3]~12_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-3]~q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add4~54\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111110000000000000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResult[-3]~12_combout\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-3]~q\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass0|Add4~54\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass0|Add4~57_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass0|Add4~58\);

-- Location: LABCELL_X18_Y64_N39
\TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-3]~12\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-3]~12_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass0|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:7:Bandpass0|Add4~57_sumout\) # (\TheRxFsk|Bandpasses:7:Bandpass0|Add4~1_sumout\) ) ) # ( 
-- !\TheRxFsk|Bandpasses:7:Bandpass0|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:7:Bandpass0|Add4~1_sumout\ & \TheRxFsk|Bandpasses:7:Bandpass0|Add4~57_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100000011000000110000001100111111001111110011111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~1_sumout\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~57_sumout\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~5_sumout\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-3]~12_combout\);

-- Location: FF_X18_Y64_N40
\TheRxFsk|Bandpasses:7:Bandpass0|Sum[-3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-3]~12_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:7:Bandpass0|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-3]~q\);

-- Location: LABCELL_X19_Y64_N39
\TheRxFsk|Bandpasses:7:Bandpass0|Add4~61\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add4~61_sumout\ = SUM(( \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-2]~DUPLICATE_q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-2]~13_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add4~58\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add4~62\ = CARRY(( \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-2]~DUPLICATE_q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-2]~13_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add4~58\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000101010101010101000000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResult[-2]~13_combout\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-2]~DUPLICATE_q\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass0|Add4~58\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass0|Add4~61_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass0|Add4~62\);

-- Location: LABCELL_X19_Y64_N57
\TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-2]~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-2]~13_combout\ = (!\TheRxFsk|Bandpasses:7:Bandpass0|Add4~1_sumout\ & (\TheRxFsk|Bandpasses:7:Bandpass0|Add4~5_sumout\ & \TheRxFsk|Bandpasses:7:Bandpass0|Add4~61_sumout\)) # 
-- (\TheRxFsk|Bandpasses:7:Bandpass0|Add4~1_sumout\ & ((\TheRxFsk|Bandpasses:7:Bandpass0|Add4~61_sumout\) # (\TheRxFsk|Bandpasses:7:Bandpass0|Add4~5_sumout\)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001011100010111000101110001011100010111000101110001011100010111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~1_sumout\,
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~5_sumout\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~61_sumout\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-2]~13_combout\);

-- Location: FF_X19_Y64_N59
\TheRxFsk|Bandpasses:7:Bandpass0|Sum[-2]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-2]~13_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:7:Bandpass0|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-2]~DUPLICATE_q\);

-- Location: LABCELL_X19_Y64_N42
\TheRxFsk|Bandpasses:7:Bandpass0|Add4~65\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add4~65_sumout\ = SUM(( \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-1]~q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-1]~14_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add4~62\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add4~66\ = CARRY(( \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-1]~q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|MultResult[-1]~14_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add4~62\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000110011001100110000000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResult[-1]~14_combout\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-1]~q\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass0|Add4~62\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass0|Add4~65_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass0|Add4~66\);

-- Location: LABCELL_X18_Y64_N45
\TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-1]~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-1]~14_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass0|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:7:Bandpass0|Add4~65_sumout\) # (\TheRxFsk|Bandpasses:7:Bandpass0|Add4~1_sumout\) ) ) # ( 
-- !\TheRxFsk|Bandpasses:7:Bandpass0|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:7:Bandpass0|Add4~1_sumout\ & \TheRxFsk|Bandpasses:7:Bandpass0|Add4~65_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100000011000000110000001100111111001111110011111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~1_sumout\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~65_sumout\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~5_sumout\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-1]~14_combout\);

-- Location: FF_X18_Y64_N46
\TheRxFsk|Bandpasses:7:Bandpass0|Sum[-1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-1]~14_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:7:Bandpass0|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-1]~q\);

-- Location: LABCELL_X19_Y64_N48
\TheRxFsk|Bandpasses:7:Bandpass0|Add4~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add4~1_sumout\ = SUM(( \TheRxFsk|Bandpasses:7:Bandpass0|Sum\(0) ) + ( !\TheRxFsk|Bandpasses:7:Bandpass0|MultResultDelayed\(0) ) + ( \TheRxFsk|Bandpasses:7:Bandpass0|Add4~6\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000001111111100000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum\(0),
	dataf => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_MultResultDelayed\(0),
	cin => \TheRxFsk|Bandpasses:7:Bandpass0|Add4~6\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass0|Add4~1_sumout\);

-- Location: LABCELL_X18_Y64_N36
\TheRxFsk|Bandpasses:7:Bandpass0|Add4~1_wirecell\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass0|Add4~1_wirecell_combout\ = !\TheRxFsk|Bandpasses:7:Bandpass0|Add4~1_sumout\

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1100110011001100110011001100110011001100110011001100110011001100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Add4~1_sumout\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass0|Add4~1_wirecell_combout\);

-- Location: FF_X18_Y64_N37
\TheRxFsk|Bandpasses:7:Bandpass0|Sum[0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass0|Add4~1_wirecell_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:7:Bandpass0|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass0|Sum\(0));

-- Location: LABCELL_X22_Y64_N27
\TheRxFsk|Mux1~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Mux1~0_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-1]~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-1]~q\ ) ) # ( !\TheRxFsk|Bandpasses:7:Bandpass0|Sum[-1]~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-1]~q\ & ( 
-- \SyncSwitchInput|Metastable\(1) ) ) ) # ( \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-1]~q\ & ( !\TheRxFsk|Bandpasses:4:Bandpass0|Sum[-1]~q\ & ( !\SyncSwitchInput|Metastable\(1) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000001111000011111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \SyncSwitchInput|ALT_INV_Metastable\(1),
	datae => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-1]~q\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-1]~q\,
	combout => \TheRxFsk|Mux1~0_combout\);

-- Location: FF_X19_Y64_N58
\TheRxFsk|Bandpasses:7:Bandpass0|Sum[-2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-2]~13_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:7:Bandpass0|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-2]~q\);

-- Location: LABCELL_X22_Y64_N6
\TheRxFsk|Mux2~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Mux2~0_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-2]~q\ & ( (!\SyncSwitchInput|Metastable\(1)) # (\TheRxFsk|Bandpasses:4:Bandpass0|Sum[-2]~q\) ) ) # ( !\TheRxFsk|Bandpasses:7:Bandpass0|Sum[-2]~q\ & ( (\SyncSwitchInput|Metastable\(1) & 
-- \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-2]~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100000011000000110000001111001111110011111100111111001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \SyncSwitchInput|ALT_INV_Metastable\(1),
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-2]~q\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-2]~q\,
	combout => \TheRxFsk|Mux2~0_combout\);

-- Location: FF_X18_Y64_N41
\TheRxFsk|Bandpasses:7:Bandpass0|Sum[-3]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-3]~12_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:7:Bandpass0|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-3]~DUPLICATE_q\);

-- Location: LABCELL_X18_Y64_N27
\TheRxFsk|Mux3~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Mux3~0_combout\ = (!\SyncSwitchInput|Metastable\(1) & (\TheRxFsk|Bandpasses:7:Bandpass0|Sum[-3]~DUPLICATE_q\)) # (\SyncSwitchInput|Metastable\(1) & ((\TheRxFsk|Bandpasses:4:Bandpass0|Sum[-3]~q\)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000101001011111000010100101111100001010010111110000101001011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \SyncSwitchInput|ALT_INV_Metastable\(1),
	datac => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-3]~DUPLICATE_q\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-3]~q\,
	combout => \TheRxFsk|Mux3~0_combout\);

-- Location: FF_X18_Y64_N17
\TheRxFsk|Bandpasses:7:Bandpass0|Sum[-4]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-4]~11_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:7:Bandpass0|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-4]~DUPLICATE_q\);

-- Location: LABCELL_X18_Y64_N24
\TheRxFsk|Mux4~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Mux4~0_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-4]~DUPLICATE_q\ & ( (!\SyncSwitchInput|Metastable\(1)) # (\TheRxFsk|Bandpasses:4:Bandpass0|Sum[-4]~q\) ) ) # ( !\TheRxFsk|Bandpasses:7:Bandpass0|Sum[-4]~DUPLICATE_q\ & ( 
-- (\SyncSwitchInput|Metastable\(1) & \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-4]~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001010101000000000101010110101010111111111010101011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \SyncSwitchInput|ALT_INV_Metastable\(1),
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-4]~q\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-4]~DUPLICATE_q\,
	combout => \TheRxFsk|Mux4~0_combout\);

-- Location: LABCELL_X23_Y64_N57
\TheRxFsk|Mux5~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Mux5~0_combout\ = (!\SyncSwitchInput|Metastable\(1) & (\TheRxFsk|Bandpasses:7:Bandpass0|Sum[-5]~q\)) # (\SyncSwitchInput|Metastable\(1) & ((\TheRxFsk|Bandpasses:4:Bandpass0|Sum[-5]~q\)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000110000111111000011000011111100001100001111110000110000111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \SyncSwitchInput|ALT_INV_Metastable\(1),
	datac => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-5]~q\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-5]~q\,
	combout => \TheRxFsk|Mux5~0_combout\);

-- Location: LABCELL_X23_Y64_N54
\TheRxFsk|Mux6~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Mux6~0_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-6]~q\ & ( (!\SyncSwitchInput|Metastable\(1)) # (\TheRxFsk|Bandpasses:4:Bandpass0|Sum[-6]~q\) ) ) # ( !\TheRxFsk|Bandpasses:7:Bandpass0|Sum[-6]~q\ & ( (\SyncSwitchInput|Metastable\(1) & 
-- \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-6]~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100000011000000110000001111001111110011111100111111001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \SyncSwitchInput|ALT_INV_Metastable\(1),
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-6]~q\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-6]~q\,
	combout => \TheRxFsk|Mux6~0_combout\);

-- Location: FF_X18_Y64_N8
\TheRxFsk|Bandpasses:7:Bandpass0|Sum[-7]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-7]~8_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:7:Bandpass0|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-7]~q\);

-- Location: LABCELL_X18_Y64_N33
\TheRxFsk|Mux7~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Mux7~0_combout\ = (!\SyncSwitchInput|Metastable\(1) & (\TheRxFsk|Bandpasses:7:Bandpass0|Sum[-7]~q\)) # (\SyncSwitchInput|Metastable\(1) & ((\TheRxFsk|Bandpasses:4:Bandpass0|Sum[-7]~q\)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000101001011111000010100101111100001010010111110000101001011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \SyncSwitchInput|ALT_INV_Metastable\(1),
	datac => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-7]~q\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-7]~q\,
	combout => \TheRxFsk|Mux7~0_combout\);

-- Location: FF_X18_Y64_N5
\TheRxFsk|Bandpasses:7:Bandpass0|Sum[-8]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass0|NextSum[-8]~7_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:7:Bandpass0|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-8]~DUPLICATE_q\);

-- Location: LABCELL_X18_Y64_N30
\TheRxFsk|Mux8~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Mux8~0_combout\ = (!\SyncSwitchInput|Metastable\(1) & (\TheRxFsk|Bandpasses:7:Bandpass0|Sum[-8]~DUPLICATE_q\)) # (\SyncSwitchInput|Metastable\(1) & ((\TheRxFsk|Bandpasses:4:Bandpass0|Sum[-8]~q\)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000101001011111000010100101111100001010010111110000101001011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \SyncSwitchInput|ALT_INV_Metastable\(1),
	datac => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-8]~DUPLICATE_q\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-8]~q\,
	combout => \TheRxFsk|Mux8~0_combout\);

-- Location: MLABCELL_X21_Y64_N6
\TheRxFsk|Mux9~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Mux9~0_combout\ = ( \SyncSwitchInput|Metastable\(1) & ( \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-9]~q\ ) ) # ( !\SyncSwitchInput|Metastable\(1) & ( \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-9]~q\ & ( \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-9]~q\ ) ) ) # 
-- ( !\SyncSwitchInput|Metastable\(1) & ( !\TheRxFsk|Bandpasses:4:Bandpass0|Sum[-9]~q\ & ( \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-9]~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001100110011000000000000000000110011001100111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-9]~q\,
	datae => \SyncSwitchInput|ALT_INV_Metastable\(1),
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-9]~q\,
	combout => \TheRxFsk|Mux9~0_combout\);

-- Location: LABCELL_X23_Y64_N48
\TheRxFsk|Mux10~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Mux10~0_combout\ = (!\SyncSwitchInput|Metastable\(1) & (\TheRxFsk|Bandpasses:7:Bandpass0|Sum[-10]~q\)) # (\SyncSwitchInput|Metastable\(1) & ((\TheRxFsk|Bandpasses:4:Bandpass0|Sum[-10]~q\)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000110000111111000011000011111100001100001111110000110000111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \SyncSwitchInput|ALT_INV_Metastable\(1),
	datac => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-10]~q\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-10]~q\,
	combout => \TheRxFsk|Mux10~0_combout\);

-- Location: LABCELL_X23_Y64_N51
\TheRxFsk|Mux11~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Mux11~0_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-11]~q\ & ( (!\SyncSwitchInput|Metastable\(1)) # (\TheRxFsk|Bandpasses:4:Bandpass0|Sum[-11]~q\) ) ) # ( !\TheRxFsk|Bandpasses:7:Bandpass0|Sum[-11]~q\ & ( (\SyncSwitchInput|Metastable\(1) 
-- & \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-11]~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100000011000000110000001111001111110011111100111111001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \SyncSwitchInput|ALT_INV_Metastable\(1),
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-11]~q\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-11]~q\,
	combout => \TheRxFsk|Mux11~0_combout\);

-- Location: LABCELL_X22_Y64_N0
\TheRxFsk|Mux12~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Mux12~0_combout\ = ( \SyncSwitchInput|Metastable\(1) & ( \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-12]~q\ ) ) # ( !\SyncSwitchInput|Metastable\(1) & ( \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-12]~q\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010101010101000011110000111101010101010101010000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-12]~q\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-12]~q\,
	datae => \SyncSwitchInput|ALT_INV_Metastable\(1),
	combout => \TheRxFsk|Mux12~0_combout\);

-- Location: LABCELL_X23_Y62_N51
\TheRxFsk|Mux13~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Mux13~0_combout\ = ( \SyncSwitchInput|Metastable\(1) & ( \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-13]~q\ ) ) # ( !\SyncSwitchInput|Metastable\(1) & ( \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-13]~q\ & ( \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-13]~q\ ) ) 
-- ) # ( !\SyncSwitchInput|Metastable\(1) & ( !\TheRxFsk|Bandpasses:4:Bandpass0|Sum[-13]~q\ & ( \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-13]~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111000000000000000000001111000011111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-13]~q\,
	datae => \SyncSwitchInput|ALT_INV_Metastable\(1),
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-13]~q\,
	combout => \TheRxFsk|Mux13~0_combout\);

-- Location: LABCELL_X22_Y64_N33
\TheRxFsk|Mux14~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Mux14~0_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-14]~q\ & ( (\TheRxFsk|Bandpasses:7:Bandpass0|Sum[-14]~q\) # (\SyncSwitchInput|Metastable\(1)) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|Sum[-14]~q\ & ( (!\SyncSwitchInput|Metastable\(1) 
-- & \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-14]~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000110000001100001111110011111100001100000011000011111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \SyncSwitchInput|ALT_INV_Metastable\(1),
	datac => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-14]~q\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-14]~q\,
	combout => \TheRxFsk|Mux14~0_combout\);

-- Location: LABCELL_X22_Y64_N12
\TheRxFsk|Mux15~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Mux15~0_combout\ = ( \SyncSwitchInput|Metastable\(1) & ( \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-15]~q\ ) ) # ( !\SyncSwitchInput|Metastable\(1) & ( \TheRxFsk|Bandpasses:4:Bandpass0|Sum[-15]~q\ & ( \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-15]~q\ ) ) 
-- ) # ( !\SyncSwitchInput|Metastable\(1) & ( !\TheRxFsk|Bandpasses:4:Bandpass0|Sum[-15]~q\ & ( \TheRxFsk|Bandpasses:7:Bandpass0|Sum[-15]~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111000000000000000000001111000011111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum[-15]~q\,
	datae => \SyncSwitchInput|ALT_INV_Metastable\(1),
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum[-15]~q\,
	combout => \TheRxFsk|Mux15~0_combout\);

-- Location: LABCELL_X23_Y64_N0
\TheRxFsk|Add0~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Add0~5_sumout\ = SUM(( !\TheRxFsk|Mux15~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:7:Bandpass0|Sum\(0)))) # (\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:4:Bandpass0|Sum\(0))))) ) + ( 
-- (!\SyncSwitchInput|Metastable\(1) & ((\TheRxFsk|Bandpasses:7:Bandpass0|Sum\(0)))) # (\SyncSwitchInput|Metastable\(1) & (\TheRxFsk|Bandpasses:4:Bandpass0|Sum\(0))) ) + ( !VCC ))
-- \TheRxFsk|Add0~6\ = CARRY(( !\TheRxFsk|Mux15~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:7:Bandpass0|Sum\(0)))) # (\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:4:Bandpass0|Sum\(0))))) ) + ( 
-- (!\SyncSwitchInput|Metastable\(1) & ((\TheRxFsk|Bandpasses:7:Bandpass0|Sum\(0)))) # (\SyncSwitchInput|Metastable\(1) & (\TheRxFsk|Bandpasses:4:Bandpass0|Sum\(0))) ) + ( !VCC ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000110010101100101000000000000000000011010111001010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum\(0),
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum\(0),
	datac => \SyncSwitchInput|ALT_INV_Metastable\(1),
	datad => \TheRxFsk|ALT_INV_Mux15~0_combout\,
	cin => GND,
	sumout => \TheRxFsk|Add0~5_sumout\,
	cout => \TheRxFsk|Add0~6\);

-- Location: LABCELL_X23_Y64_N3
\TheRxFsk|Add0~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Add0~9_sumout\ = SUM(( !\TheRxFsk|Mux14~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:7:Bandpass0|Sum\(0)))) # (\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:4:Bandpass0|Sum\(0))))) ) + ( GND ) + ( 
-- \TheRxFsk|Add0~6\ ))
-- \TheRxFsk|Add0~10\ = CARRY(( !\TheRxFsk|Mux14~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:7:Bandpass0|Sum\(0)))) # (\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:4:Bandpass0|Sum\(0))))) ) + ( GND ) + ( 
-- \TheRxFsk|Add0~6\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000011010111001010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum\(0),
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum\(0),
	datac => \SyncSwitchInput|ALT_INV_Metastable\(1),
	datad => \TheRxFsk|ALT_INV_Mux14~0_combout\,
	cin => \TheRxFsk|Add0~6\,
	sumout => \TheRxFsk|Add0~9_sumout\,
	cout => \TheRxFsk|Add0~10\);

-- Location: LABCELL_X23_Y64_N6
\TheRxFsk|Add0~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Add0~13_sumout\ = SUM(( !\TheRxFsk|Mux13~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:7:Bandpass0|Sum\(0)))) # (\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:4:Bandpass0|Sum\(0))))) ) + ( GND ) + ( 
-- \TheRxFsk|Add0~10\ ))
-- \TheRxFsk|Add0~14\ = CARRY(( !\TheRxFsk|Mux13~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:7:Bandpass0|Sum\(0)))) # (\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:4:Bandpass0|Sum\(0))))) ) + ( GND ) + ( 
-- \TheRxFsk|Add0~10\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000011010111001010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum\(0),
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum\(0),
	datac => \SyncSwitchInput|ALT_INV_Metastable\(1),
	datad => \TheRxFsk|ALT_INV_Mux13~0_combout\,
	cin => \TheRxFsk|Add0~10\,
	sumout => \TheRxFsk|Add0~13_sumout\,
	cout => \TheRxFsk|Add0~14\);

-- Location: LABCELL_X23_Y64_N9
\TheRxFsk|Add0~17\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Add0~17_sumout\ = SUM(( GND ) + ( !\TheRxFsk|Mux12~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:7:Bandpass0|Sum\(0)))) # (\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:4:Bandpass0|Sum\(0))))) ) + ( 
-- \TheRxFsk|Add0~14\ ))
-- \TheRxFsk|Add0~18\ = CARRY(( GND ) + ( !\TheRxFsk|Mux12~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:7:Bandpass0|Sum\(0)))) # (\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:4:Bandpass0|Sum\(0))))) ) + ( 
-- \TheRxFsk|Add0~14\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000110010100011010100000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum\(0),
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum\(0),
	datac => \SyncSwitchInput|ALT_INV_Metastable\(1),
	dataf => \TheRxFsk|ALT_INV_Mux12~0_combout\,
	cin => \TheRxFsk|Add0~14\,
	sumout => \TheRxFsk|Add0~17_sumout\,
	cout => \TheRxFsk|Add0~18\);

-- Location: LABCELL_X23_Y64_N12
\TheRxFsk|Add0~21\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Add0~21_sumout\ = SUM(( GND ) + ( !\TheRxFsk|Mux11~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:7:Bandpass0|Sum\(0)))) # (\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:4:Bandpass0|Sum\(0))))) ) + ( 
-- \TheRxFsk|Add0~18\ ))
-- \TheRxFsk|Add0~22\ = CARRY(( GND ) + ( !\TheRxFsk|Mux11~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:7:Bandpass0|Sum\(0)))) # (\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:4:Bandpass0|Sum\(0))))) ) + ( 
-- \TheRxFsk|Add0~18\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000110010100011010100000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum\(0),
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum\(0),
	datac => \SyncSwitchInput|ALT_INV_Metastable\(1),
	dataf => \TheRxFsk|ALT_INV_Mux11~0_combout\,
	cin => \TheRxFsk|Add0~18\,
	sumout => \TheRxFsk|Add0~21_sumout\,
	cout => \TheRxFsk|Add0~22\);

-- Location: LABCELL_X23_Y64_N15
\TheRxFsk|Add0~25\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Add0~25_sumout\ = SUM(( GND ) + ( !\TheRxFsk|Mux10~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:7:Bandpass0|Sum\(0)))) # (\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:4:Bandpass0|Sum\(0))))) ) + ( 
-- \TheRxFsk|Add0~22\ ))
-- \TheRxFsk|Add0~26\ = CARRY(( GND ) + ( !\TheRxFsk|Mux10~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:7:Bandpass0|Sum\(0)))) # (\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:4:Bandpass0|Sum\(0))))) ) + ( 
-- \TheRxFsk|Add0~22\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000110010100011010100000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum\(0),
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum\(0),
	datac => \SyncSwitchInput|ALT_INV_Metastable\(1),
	dataf => \TheRxFsk|ALT_INV_Mux10~0_combout\,
	cin => \TheRxFsk|Add0~22\,
	sumout => \TheRxFsk|Add0~25_sumout\,
	cout => \TheRxFsk|Add0~26\);

-- Location: LABCELL_X23_Y64_N18
\TheRxFsk|Add0~29\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Add0~29_sumout\ = SUM(( !\TheRxFsk|Mux9~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:7:Bandpass0|Sum\(0)))) # (\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:4:Bandpass0|Sum\(0))))) ) + ( GND ) + ( 
-- \TheRxFsk|Add0~26\ ))
-- \TheRxFsk|Add0~30\ = CARRY(( !\TheRxFsk|Mux9~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:7:Bandpass0|Sum\(0)))) # (\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:4:Bandpass0|Sum\(0))))) ) + ( GND ) + ( 
-- \TheRxFsk|Add0~26\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000011010111001010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum\(0),
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum\(0),
	datac => \SyncSwitchInput|ALT_INV_Metastable\(1),
	datad => \TheRxFsk|ALT_INV_Mux9~0_combout\,
	cin => \TheRxFsk|Add0~26\,
	sumout => \TheRxFsk|Add0~29_sumout\,
	cout => \TheRxFsk|Add0~30\);

-- Location: LABCELL_X23_Y64_N21
\TheRxFsk|Add0~33\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Add0~33_sumout\ = SUM(( !\TheRxFsk|Mux8~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:7:Bandpass0|Sum\(0)))) # (\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:4:Bandpass0|Sum\(0))))) ) + ( GND ) + ( 
-- \TheRxFsk|Add0~30\ ))
-- \TheRxFsk|Add0~34\ = CARRY(( !\TheRxFsk|Mux8~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:7:Bandpass0|Sum\(0)))) # (\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:4:Bandpass0|Sum\(0))))) ) + ( GND ) + ( 
-- \TheRxFsk|Add0~30\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000011010111001010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum\(0),
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum\(0),
	datac => \SyncSwitchInput|ALT_INV_Metastable\(1),
	datad => \TheRxFsk|ALT_INV_Mux8~0_combout\,
	cin => \TheRxFsk|Add0~30\,
	sumout => \TheRxFsk|Add0~33_sumout\,
	cout => \TheRxFsk|Add0~34\);

-- Location: LABCELL_X23_Y64_N24
\TheRxFsk|Add0~37\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Add0~37_sumout\ = SUM(( GND ) + ( !\TheRxFsk|Mux7~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:7:Bandpass0|Sum\(0)))) # (\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:4:Bandpass0|Sum\(0))))) ) + ( 
-- \TheRxFsk|Add0~34\ ))
-- \TheRxFsk|Add0~38\ = CARRY(( GND ) + ( !\TheRxFsk|Mux7~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:7:Bandpass0|Sum\(0)))) # (\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:4:Bandpass0|Sum\(0))))) ) + ( 
-- \TheRxFsk|Add0~34\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000110010100011010100000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum\(0),
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum\(0),
	datac => \SyncSwitchInput|ALT_INV_Metastable\(1),
	dataf => \TheRxFsk|ALT_INV_Mux7~0_combout\,
	cin => \TheRxFsk|Add0~34\,
	sumout => \TheRxFsk|Add0~37_sumout\,
	cout => \TheRxFsk|Add0~38\);

-- Location: LABCELL_X23_Y64_N27
\TheRxFsk|Add0~41\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Add0~41_sumout\ = SUM(( !\TheRxFsk|Mux6~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:7:Bandpass0|Sum\(0)))) # (\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:4:Bandpass0|Sum\(0))))) ) + ( GND ) + ( 
-- \TheRxFsk|Add0~38\ ))
-- \TheRxFsk|Add0~42\ = CARRY(( !\TheRxFsk|Mux6~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:7:Bandpass0|Sum\(0)))) # (\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:4:Bandpass0|Sum\(0))))) ) + ( GND ) + ( 
-- \TheRxFsk|Add0~38\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000011010111001010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum\(0),
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum\(0),
	datac => \SyncSwitchInput|ALT_INV_Metastable\(1),
	datad => \TheRxFsk|ALT_INV_Mux6~0_combout\,
	cin => \TheRxFsk|Add0~38\,
	sumout => \TheRxFsk|Add0~41_sumout\,
	cout => \TheRxFsk|Add0~42\);

-- Location: LABCELL_X23_Y64_N30
\TheRxFsk|Add0~45\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Add0~45_sumout\ = SUM(( !\TheRxFsk|Mux5~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:7:Bandpass0|Sum\(0)))) # (\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:4:Bandpass0|Sum\(0))))) ) + ( GND ) + ( 
-- \TheRxFsk|Add0~42\ ))
-- \TheRxFsk|Add0~46\ = CARRY(( !\TheRxFsk|Mux5~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:7:Bandpass0|Sum\(0)))) # (\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:4:Bandpass0|Sum\(0))))) ) + ( GND ) + ( 
-- \TheRxFsk|Add0~42\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000011010111001010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum\(0),
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum\(0),
	datac => \SyncSwitchInput|ALT_INV_Metastable\(1),
	datad => \TheRxFsk|ALT_INV_Mux5~0_combout\,
	cin => \TheRxFsk|Add0~42\,
	sumout => \TheRxFsk|Add0~45_sumout\,
	cout => \TheRxFsk|Add0~46\);

-- Location: LABCELL_X23_Y64_N33
\TheRxFsk|Add0~49\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Add0~49_sumout\ = SUM(( !\TheRxFsk|Mux4~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:7:Bandpass0|Sum\(0)))) # (\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:4:Bandpass0|Sum\(0))))) ) + ( GND ) + ( 
-- \TheRxFsk|Add0~46\ ))
-- \TheRxFsk|Add0~50\ = CARRY(( !\TheRxFsk|Mux4~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:7:Bandpass0|Sum\(0)))) # (\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:4:Bandpass0|Sum\(0))))) ) + ( GND ) + ( 
-- \TheRxFsk|Add0~46\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000011010111001010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum\(0),
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum\(0),
	datac => \SyncSwitchInput|ALT_INV_Metastable\(1),
	datad => \TheRxFsk|ALT_INV_Mux4~0_combout\,
	cin => \TheRxFsk|Add0~46\,
	sumout => \TheRxFsk|Add0~49_sumout\,
	cout => \TheRxFsk|Add0~50\);

-- Location: LABCELL_X23_Y64_N36
\TheRxFsk|Add0~53\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Add0~53_sumout\ = SUM(( !\TheRxFsk|Mux3~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:7:Bandpass0|Sum\(0)))) # (\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:4:Bandpass0|Sum\(0))))) ) + ( GND ) + ( 
-- \TheRxFsk|Add0~50\ ))
-- \TheRxFsk|Add0~54\ = CARRY(( !\TheRxFsk|Mux3~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:7:Bandpass0|Sum\(0)))) # (\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:4:Bandpass0|Sum\(0))))) ) + ( GND ) + ( 
-- \TheRxFsk|Add0~50\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000011010111001010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum\(0),
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum\(0),
	datac => \SyncSwitchInput|ALT_INV_Metastable\(1),
	datad => \TheRxFsk|ALT_INV_Mux3~0_combout\,
	cin => \TheRxFsk|Add0~50\,
	sumout => \TheRxFsk|Add0~53_sumout\,
	cout => \TheRxFsk|Add0~54\);

-- Location: LABCELL_X23_Y64_N39
\TheRxFsk|Add0~57\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Add0~57_sumout\ = SUM(( !\TheRxFsk|Mux2~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:7:Bandpass0|Sum\(0)))) # (\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:4:Bandpass0|Sum\(0))))) ) + ( GND ) + ( 
-- \TheRxFsk|Add0~54\ ))
-- \TheRxFsk|Add0~58\ = CARRY(( !\TheRxFsk|Mux2~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:7:Bandpass0|Sum\(0)))) # (\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:4:Bandpass0|Sum\(0))))) ) + ( GND ) + ( 
-- \TheRxFsk|Add0~54\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000011010111001010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum\(0),
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum\(0),
	datac => \SyncSwitchInput|ALT_INV_Metastable\(1),
	datad => \TheRxFsk|ALT_INV_Mux2~0_combout\,
	cin => \TheRxFsk|Add0~54\,
	sumout => \TheRxFsk|Add0~57_sumout\,
	cout => \TheRxFsk|Add0~58\);

-- Location: LABCELL_X23_Y64_N42
\TheRxFsk|Add0~61\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Add0~61_sumout\ = SUM(( !\TheRxFsk|Mux1~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:7:Bandpass0|Sum\(0)))) # (\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:4:Bandpass0|Sum\(0))))) ) + ( GND ) + ( 
-- \TheRxFsk|Add0~58\ ))
-- \TheRxFsk|Add0~62\ = CARRY(( !\TheRxFsk|Mux1~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:7:Bandpass0|Sum\(0)))) # (\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:4:Bandpass0|Sum\(0))))) ) + ( GND ) + ( 
-- \TheRxFsk|Add0~58\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000011010111001010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_Sum\(0),
	datab => \TheRxFsk|Bandpasses:7:Bandpass0|ALT_INV_Sum\(0),
	datac => \SyncSwitchInput|ALT_INV_Metastable\(1),
	datad => \TheRxFsk|ALT_INV_Mux1~0_combout\,
	cin => \TheRxFsk|Add0~58\,
	sumout => \TheRxFsk|Add0~61_sumout\,
	cout => \TheRxFsk|Add0~62\);

-- Location: LABCELL_X23_Y64_N45
\TheRxFsk|Add0~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Add0~1_sumout\ = SUM(( GND ) + ( GND ) + ( \TheRxFsk|Add0~62\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	cin => \TheRxFsk|Add0~62\,
	sumout => \TheRxFsk|Add0~1_sumout\);

-- Location: M10K_X26_Y61_N0
\TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a0\ : cyclonev_ram_block
-- pragma translate_off
GENERIC MAP (
	mem_init4 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	mem_init3 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	mem_init2 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000039BFFD8A0004F00144FFF94FFE8300165000FEFFDF1FFFF30025AFFEE8FFE0B002400010EFFCE30006C0033CFFDF6FFD920038E000E0FFBA70013F00418FFC9EFFD410051B00068FFA450027C004F4FFAEFFFD49006E9FFF72FF8E70042D00582FF8DAFFDCA008DEFFE07FF7A60065B005BBFF67DFFEC800AC3FFC02FF6A2008E30",
	mem_init1 => "0569FF3F80005600C8DFF975FF62B00BDF00473FF17F0029100DFEFF66DFF63A00EEC002DAFEF2B0056F00ED9FF30FFF70B011E500076FED4C008C000F04FEF83FF8A0014A8FFD60FEC0400C8C00E6EFEC09FFB1A016FDFF9DBFEB950106900CD7FE8E1FFE3701885FF5D7FEC020143A00A73FE64D001FF0193BFF1BAFED68017A80074AFE47D00610018F0FEDA3FEFC401A830037AFE39100A60017AAFEA0DFF2EE01C81FFF41FE3BD00E8E01560FE708FF6B901D98FFAF0FE4DF0124501245FE4DFFFAF001D98FF6B9FE7080156000E8EFE3BDFFF4101C81FF2EEFEA0D017AA00A60FE3910037A01A83FEFC4FEDA3018F000610FE47D0074A017A8FED68FF1",
	mem_init0 => "BA0193B001FFFE64D00A730143AFEC02FF5D701885FFE37FE8E100CD701069FEB95FF9DB016FDFFB1AFEC0900E6E00C8CFEC04FFD60014A8FF8A0FEF8300F04008C0FED4C00076011E5FF70BFF30F00ED90056FFEF2B002DA00EECFF63AFF66D00DFE00291FF17F0047300BDFFF62BFF97500C8D00056FF3F800569008E3FF6A2FFC0200AC3FFEC8FF67D005BB0065BFF7A6FFE07008DEFFDCAFF8DA005820042DFF8E7FFF72006E9FFD49FFAEF004F40027CFFA45000680051BFFD41FFC9E004180013FFFBA7000E00038EFFD92FFDF60033C0006CFFCE30010E00240FFE0BFFEE80025AFFFF3FFDF1000FE00165FFE83FFF94001440004FFFD8A0039B00200",
	data_interleave_offset_in_bits => 1,
	data_interleave_width_in_bits => 1,
	init_file => "db/TbdRxFskBasic.ram1_DspFir_2df41c30.hdl.mif",
	init_file_layout => "port_a",
	logical_ram_name => "RxFsk:TheRxFsk|DspFir:\Bandpasses:4:Bandpass1|altsyncram:CoefMemory_rtl_0|altsyncram_2nd1:auto_generated|ALTSYNCRAM",
	operation_mode => "rom",
	port_a_address_clear => "none",
	port_a_address_width => 9,
	port_a_byte_enable_clock => "none",
	port_a_data_out_clear => "none",
	port_a_data_out_clock => "none",
	port_a_data_width => 20,
	port_a_first_address => 0,
	port_a_first_bit_number => 0,
	port_a_last_address => 511,
	port_a_logical_ram_depth => 258,
	port_a_logical_ram_width => 16,
	port_a_read_during_write_mode => "new_data_no_nbe_read",
	port_a_write_enable_clock => "none",
	port_b_address_width => 9,
	port_b_data_width => 20,
	ram_block_type => "M20K")
-- pragma translate_on
PORT MAP (
	portare => VCC,
	clk0 => \iClk~inputCLKENA0_outclk\,
	portaaddr => \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a0_PORTAADDR_bus\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	portadataout => \TheRxFsk|Bandpasses:4:Bandpass1|CoefMemory_rtl_0|auto_generated|ram_block1a0_PORTADATAOUT_bus\);

-- Location: M10K_X14_Y63_N0
\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a0\ : cyclonev_ram_block
-- pragma translate_off
GENERIC MAP (
	mem_init4 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	mem_init3 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	mem_init2 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	mem_init1 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	mem_init0 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	data_interleave_offset_in_bits => 1,
	data_interleave_width_in_bits => 1,
	init_file => "db/TbdRxFskBasic.ram0_DspFir_2df41c30.hdl.mif",
	init_file_layout => "port_a",
	logical_ram_name => "RxFsk:TheRxFsk|DspFir:\Bandpasses:4:Bandpass1|altsyncram:SampleMemory_rtl_0|altsyncram_cbs1:auto_generated|ALTSYNCRAM",
	mixed_port_feed_through_mode => "old",
	operation_mode => "dual_port",
	port_a_address_clear => "none",
	port_a_address_width => 9,
	port_a_byte_enable_clock => "none",
	port_a_data_out_clear => "none",
	port_a_data_out_clock => "none",
	port_a_data_width => 20,
	port_a_first_address => 0,
	port_a_first_bit_number => 0,
	port_a_last_address => 511,
	port_a_logical_ram_depth => 258,
	port_a_logical_ram_width => 16,
	port_a_read_during_write_mode => "new_data_no_nbe_read",
	port_b_address_clear => "none",
	port_b_address_clock => "clock0",
	port_b_address_width => 9,
	port_b_data_out_clear => "none",
	port_b_data_out_clock => "none",
	port_b_data_width => 20,
	port_b_first_address => 0,
	port_b_first_bit_number => 0,
	port_b_last_address => 511,
	port_b_logical_ram_depth => 258,
	port_b_logical_ram_width => 16,
	port_b_read_during_write_mode => "new_data_no_nbe_read",
	port_b_read_enable_clock => "clock0",
	ram_block_type => "M20K")
-- pragma translate_on
PORT MAP (
	portawe => \TheI2sToPar|ValL~q\,
	portbre => VCC,
	clk0 => \iClk~inputCLKENA0_outclk\,
	portadatain => \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTADATAIN_bus\,
	portaaddr => \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTAADDR_bus\,
	portbaddr => \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBADDR_bus\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	portbdataout => \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\);

-- Location: LABCELL_X16_Y62_N51
\TheRxFsk|Bandpasses:4:Bandpass1|Sample[-15]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-15]~0_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a0~portbdataout\ ) ) # ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a0~portbdataout\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-15]~q\ ) ) ) # ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( !\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a0~portbdataout\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-15]~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010101010101000000000000000001010101010101011111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-15]~q\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a0~portbdataout\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-15]~0_combout\);

-- Location: LABCELL_X18_Y63_N3
\TheRxFsk|Bandpasses:4:Bandpass1|Sample[-14]~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-14]~1_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a1\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-14]~q\ ) ) # ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a1\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-14]~q\ & ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ ) ) ) # ( 
-- \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a1\ & ( !\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-14]~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000010101010101010110101010101010101111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a1\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-14]~q\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-14]~1_combout\);

-- Location: LABCELL_X19_Y63_N6
\TheRxFsk|Bandpasses:4:Bandpass1|Sample[-13]~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-13]~2_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-13]~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a2\ ) ) 
-- ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-13]~q\ ) ) # ( \TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( !\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-13]~q\ & ( 
-- \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a2\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000011110000111111111111111111110000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a2\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-13]~q\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-13]~2_combout\);

-- Location: LABCELL_X18_Y61_N6
\TheRxFsk|Bandpasses:4:Bandpass1|Sample[-12]~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-12]~3_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-12]~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a3\ ) ) 
-- ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-12]~q\ ) ) # ( \TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( !\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-12]~q\ & ( 
-- \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a3\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000011110000111111111111111111110000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a3\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-12]~q\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-12]~3_combout\);

-- Location: MLABCELL_X15_Y63_N12
\TheRxFsk|Bandpasses:4:Bandpass1|Sample[-11]~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-11]~4_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a4~portbdataout\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-11]~q\) # 
-- (\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a4~portbdataout\ & ( (!\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & 
-- \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-11]~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000110000001100000011000000110000111111001111110011111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-11]~q\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a4~portbdataout\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-11]~4_combout\);

-- Location: LABCELL_X19_Y62_N6
\TheRxFsk|Bandpasses:4:Bandpass1|Sample[-10]~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-10]~5_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a5\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-10]~q\ ) ) # ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a5\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-10]~q\ & ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ ) ) ) # ( 
-- \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a5\ & ( !\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-10]~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000001100110011001111001100110011001111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a5\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-10]~q\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-10]~5_combout\);

-- Location: LABCELL_X18_Y63_N54
\TheRxFsk|Bandpasses:4:Bandpass1|Sample[-9]~6\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-9]~6_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a6\ ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & 
-- ( \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a6\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-9]~q\ ) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a6\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-9]~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111000000000000000000001111000011111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-9]~q\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a6\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-9]~6_combout\);

-- Location: LABCELL_X18_Y62_N9
\TheRxFsk|Bandpasses:4:Bandpass1|Sample[-8]~7\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-8]~7_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a7\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-8]~q\ ) ) # ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a7\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-8]~q\ & ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ ) ) ) # ( 
-- \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a7\ & ( !\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-8]~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000011110000111111110000111100001111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a7\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-8]~q\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-8]~7_combout\);

-- Location: LABCELL_X17_Y63_N21
\TheRxFsk|Bandpasses:4:Bandpass1|Sample[-7]~8\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-7]~8_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a8\ ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & 
-- ( \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a8\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-7]~q\ ) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a8\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-7]~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111000000000000000000001111000011111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-7]~q\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a8\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-7]~8_combout\);

-- Location: LABCELL_X16_Y61_N24
\TheRxFsk|Bandpasses:4:Bandpass1|Sample[-6]~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-6]~9_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-6]~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a9\ ) ) # ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-6]~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a9\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ ) ) ) # ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-6]~q\ & 
-- ( !\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a9\ & ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000110011001100110000110011001100111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-6]~q\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a9\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-6]~9_combout\);

-- Location: LABCELL_X18_Y63_N24
\TheRxFsk|Bandpasses:4:Bandpass1|Sample[-5]~10\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-5]~10_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a10\ ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ 
-- & ( \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a10\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-5]~q\ ) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a10\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-5]~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111000000000000000000001111000011111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-5]~q\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a10\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-5]~10_combout\);

-- Location: MLABCELL_X15_Y63_N18
\TheRxFsk|Bandpasses:4:Bandpass1|Sample[-4]~11\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-4]~11_combout\ = (!\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ((\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-4]~q\))) # (\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & 
-- (\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a11\))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001101100011011000110110001101100011011000110110001101100011011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	datab => \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a11\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-4]~q\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-4]~11_combout\);

-- Location: LABCELL_X17_Y65_N24
\TheRxFsk|Bandpasses:4:Bandpass1|Sample[-3]~12\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-3]~12_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a12\ ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ 
-- & ( \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a12\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-3]~q\ ) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a12\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-3]~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111000000000000000000001111000011111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-3]~q\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a12\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-3]~12_combout\);

-- Location: LABCELL_X19_Y63_N51
\TheRxFsk|Bandpasses:4:Bandpass1|Sample[-2]~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-2]~13_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a13\ ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ 
-- & ( \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a13\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-2]~q\ ) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a13\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-2]~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010101010101000000000000000001010101010101011111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-2]~q\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a13\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-2]~13_combout\);

-- Location: LABCELL_X19_Y63_N42
\TheRxFsk|Bandpasses:4:Bandpass1|Sample[-1]~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-1]~14_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a14\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\) # (\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-1]~q\) ) 
-- ) # ( !\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a14\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-1]~q\ & !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011000000110000001100000011000000111111001111110011111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-1]~q\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a14\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|Sample[-1]~14_combout\);

-- Location: MLABCELL_X15_Y62_N9
\TheRxFsk|Bandpasses:4:Bandpass1|Sample[0]~15\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Sample[0]~15_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[0]~DUPLICATE_q\ & ( (!\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\) # 
-- (\TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a15\) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[0]~DUPLICATE_q\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & 
-- \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a15\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100000011000000110000001111001111110011111100111111001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a15\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[0]~DUPLICATE_q\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|Sample[0]~15_combout\);

-- Location: DSP_X20_Y59_N0
\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8\ : cyclonev_mac
-- pragma translate_off
GENERIC MAP (
	accumulate_clock => "none",
	ax_clock => "none",
	ax_width => 18,
	ay_scan_in_clock => "none",
	ay_scan_in_width => 19,
	ay_use_scan_in => "false",
	az_clock => "none",
	bx_clock => "none",
	by_clock => "none",
	by_use_scan_in => "false",
	bz_clock => "none",
	coef_a_0 => 0,
	coef_a_1 => 0,
	coef_a_2 => 0,
	coef_a_3 => 0,
	coef_a_4 => 0,
	coef_a_5 => 0,
	coef_a_6 => 0,
	coef_a_7 => 0,
	coef_b_0 => 0,
	coef_b_1 => 0,
	coef_b_2 => 0,
	coef_b_3 => 0,
	coef_b_4 => 0,
	coef_b_5 => 0,
	coef_b_6 => 0,
	coef_b_7 => 0,
	coef_sel_a_clock => "none",
	coef_sel_b_clock => "none",
	delay_scan_out_ay => "false",
	delay_scan_out_by => "false",
	enable_double_accum => "false",
	load_const_clock => "none",
	load_const_value => 0,
	mode_sub_location => 0,
	negate_clock => "none",
	operand_source_max => "input",
	operand_source_may => "input",
	operand_source_mbx => "input",
	operand_source_mby => "input",
	operation_mode => "m18x18_full",
	output_clock => "none",
	preadder_subtract_a => "false",
	preadder_subtract_b => "false",
	result_a_width => 64,
	signed_max => "true",
	signed_may => "true",
	signed_mbx => "false",
	signed_mby => "false",
	sub_clock => "none",
	use_chainadder => "false")
-- pragma translate_on
PORT MAP (
	sub => GND,
	negate => GND,
	ax => \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_AX_bus\,
	ay => \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_AY_bus\,
	resulta => \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_RESULTA_bus\);

-- Location: MLABCELL_X21_Y59_N45
\TheRxFsk|Bandpasses:4:Bandpass1|vAdd~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|vAdd~2_combout\ = ( !\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~12\ & ( !\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~8_resulta\ & ( (!\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~21\ & (!\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~10\ & 
-- !\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~11\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1000000010000000000000000000000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~21\,
	datab => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~10\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~11\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~12\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~8_resulta\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|vAdd~2_combout\);

-- Location: MLABCELL_X21_Y59_N0
\TheRxFsk|Bandpasses:4:Bandpass1|vAdd~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|vAdd~1_combout\ = ( !\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~14\ & ( !\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~9\ & ( (!\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~15\ & (!\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~18\ & 
-- (!\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~17\ & !\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~16\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1000000000000000000000000000000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~15\,
	datab => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~18\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~17\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~16\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~14\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~9\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|vAdd~1_combout\);

-- Location: LABCELL_X19_Y59_N54
\TheRxFsk|Bandpasses:4:Bandpass1|vAdd~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|vAdd~0_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass1|vAdd~2_combout\ & ( \TheRxFsk|Bandpasses:4:Bandpass1|vAdd~1_combout\ & ( (((\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~19\) # (\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~13\)) # 
-- (\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~22\)) # (\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~20\) ) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass1|vAdd~2_combout\ & ( \TheRxFsk|Bandpasses:4:Bandpass1|vAdd~1_combout\ ) ) # ( 
-- \TheRxFsk|Bandpasses:4:Bandpass1|vAdd~2_combout\ & ( !\TheRxFsk|Bandpasses:4:Bandpass1|vAdd~1_combout\ ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass1|vAdd~2_combout\ & ( !\TheRxFsk|Bandpasses:4:Bandpass1|vAdd~1_combout\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111111111111111111111111111111111111111111110111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~20\,
	datab => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~22\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~13\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~19\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_vAdd~2_combout\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_vAdd~1_combout\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|vAdd~0_combout\);

-- Location: LABCELL_X19_Y59_N0
\TheRxFsk|Bandpasses:4:Bandpass1|Add3~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add3~13_sumout\ = SUM(( (\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~39\ & \TheRxFsk|Bandpasses:4:Bandpass1|vAdd~0_combout\) ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~23\ ) + ( !VCC ))
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add3~14\ = CARRY(( (\TheRxFsk|Bandpasses:4:Bandpass1|Mult0~39\ & \TheRxFsk|Bandpasses:4:Bandpass1|vAdd~0_combout\) ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~23\ ) + ( !VCC ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~39\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~23\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_vAdd~0_combout\,
	cin => GND,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~13_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~14\);

-- Location: LABCELL_X19_Y59_N3
\TheRxFsk|Bandpasses:4:Bandpass1|Add3~17\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add3~17_sumout\ = SUM(( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~24\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add3~14\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add3~18\ = CARRY(( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~24\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add3~14\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~24\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~14\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~17_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~18\);

-- Location: LABCELL_X19_Y59_N6
\TheRxFsk|Bandpasses:4:Bandpass1|Add3~21\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add3~21_sumout\ = SUM(( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~25\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add3~18\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add3~22\ = CARRY(( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~25\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add3~18\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~25\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~18\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~21_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~22\);

-- Location: LABCELL_X19_Y59_N9
\TheRxFsk|Bandpasses:4:Bandpass1|Add3~25\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add3~25_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~26\ ) + ( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add3~22\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add3~26\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~26\ ) + ( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add3~22\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~26\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~22\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~25_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~26\);

-- Location: LABCELL_X19_Y59_N12
\TheRxFsk|Bandpasses:4:Bandpass1|Add3~29\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add3~29_sumout\ = SUM(( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~27\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add3~26\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add3~30\ = CARRY(( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~27\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add3~26\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~27\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~26\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~29_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~30\);

-- Location: LABCELL_X19_Y59_N15
\TheRxFsk|Bandpasses:4:Bandpass1|Add3~33\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add3~33_sumout\ = SUM(( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~28\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add3~30\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add3~34\ = CARRY(( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~28\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add3~30\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~28\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~30\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~33_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~34\);

-- Location: LABCELL_X19_Y59_N18
\TheRxFsk|Bandpasses:4:Bandpass1|Add3~37\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add3~37_sumout\ = SUM(( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~29\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add3~34\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add3~38\ = CARRY(( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~29\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add3~34\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~29\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~34\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~37_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~38\);

-- Location: LABCELL_X19_Y59_N21
\TheRxFsk|Bandpasses:4:Bandpass1|Add3~41\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add3~41_sumout\ = SUM(( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~30\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add3~38\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add3~42\ = CARRY(( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~30\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add3~38\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~30\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~38\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~41_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~42\);

-- Location: LABCELL_X19_Y59_N24
\TheRxFsk|Bandpasses:4:Bandpass1|Add3~45\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add3~45_sumout\ = SUM(( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~31\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add3~42\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add3~46\ = CARRY(( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~31\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add3~42\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~31\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~42\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~45_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~46\);

-- Location: LABCELL_X19_Y59_N27
\TheRxFsk|Bandpasses:4:Bandpass1|Add3~49\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add3~49_sumout\ = SUM(( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~32\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add3~46\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add3~50\ = CARRY(( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~32\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add3~46\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~32\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~46\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~49_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~50\);

-- Location: LABCELL_X19_Y59_N30
\TheRxFsk|Bandpasses:4:Bandpass1|Add3~53\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add3~53_sumout\ = SUM(( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~33\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add3~50\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add3~54\ = CARRY(( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~33\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add3~50\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~33\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~50\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~53_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~54\);

-- Location: LABCELL_X19_Y59_N33
\TheRxFsk|Bandpasses:4:Bandpass1|Add3~57\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add3~57_sumout\ = SUM(( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~34\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add3~54\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add3~58\ = CARRY(( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~34\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add3~54\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~34\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~54\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~57_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~58\);

-- Location: LABCELL_X19_Y59_N36
\TheRxFsk|Bandpasses:4:Bandpass1|Add3~61\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add3~61_sumout\ = SUM(( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~35\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add3~58\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add3~62\ = CARRY(( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~35\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add3~58\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~35\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~58\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~61_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~62\);

-- Location: LABCELL_X19_Y59_N39
\TheRxFsk|Bandpasses:4:Bandpass1|Add3~65\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add3~65_sumout\ = SUM(( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~36\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add3~62\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add3~66\ = CARRY(( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~36\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add3~62\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000101010101010101000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~36\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~62\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~65_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~66\);

-- Location: LABCELL_X19_Y59_N42
\TheRxFsk|Bandpasses:4:Bandpass1|Add3~69\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add3~69_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~37\ ) + ( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add3~66\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add3~70\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~37\ ) + ( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add3~66\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~37\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~66\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~69_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~70\);

-- Location: LABCELL_X19_Y59_N45
\TheRxFsk|Bandpasses:4:Bandpass1|Add3~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add3~9_sumout\ = SUM(( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~38\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add3~70\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add3~10\ = CARRY(( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~38\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add3~70\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000101010101010101000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~38\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~70\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~9_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~10\);

-- Location: LABCELL_X19_Y59_N48
\TheRxFsk|Bandpasses:4:Bandpass1|Add3~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add3~5_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~39\ ) + ( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add3~10\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add3~6\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~39\ ) + ( GND ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add3~10\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~39\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~10\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~5_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~6\);

-- Location: LABCELL_X19_Y59_N51
\TheRxFsk|Bandpasses:4:Bandpass1|Add3~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add3~1_sumout\ = SUM(( VCC ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Mult0~39\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add3~6\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000001111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Mult0~39\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~6\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~1_sumout\);

-- Location: LABCELL_X22_Y59_N0
\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[0]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[0]~0_combout\ = ( !\TheRxFsk|Bandpasses:4:Bandpass1|Add3~1_sumout\ )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111111111111111111111111111100000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add3~1_sumout\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[0]~0_combout\);

-- Location: FF_X22_Y59_N1
\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[0]~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed\(0));

-- Location: FF_X19_Y59_N46
\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_NEW_REG84\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~9_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM85\);

-- Location: FF_X19_Y59_N53
\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_NEW_REG80\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~1_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM81\);

-- Location: FF_X19_Y59_N49
\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_NEW_REG82\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~5_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM83\);

-- Location: FF_X19_Y59_N43
\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-1]_NEW_REG100\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~69_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-1]_OTERM101\);

-- Location: LABCELL_X19_Y60_N18
\TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-1]~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-1]~14_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM83\ & ( \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-1]_OTERM101\ & ( 
-- (\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM81\) # (\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM85\) ) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM83\ & ( 
-- \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-1]_OTERM101\ & ( \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM81\ ) ) ) # ( \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM83\ & ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-1]_OTERM101\ & ( \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM81\ ) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM83\ & ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-1]_OTERM101\ & ( (\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM85\ & \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM81\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100000011000011110000111100001111000011110011111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM85\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM81\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM83\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-1]_OTERM101\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-1]~14_combout\);

-- Location: FF_X19_Y59_N40
\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-2]_NEW_REG106\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~65_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-2]_OTERM107\);

-- Location: LABCELL_X19_Y60_N39
\TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-2]~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-2]~13_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-2]_OTERM107\ & ( ((\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM83\ & 
-- \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM85\)) # (\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM81\) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-2]_OTERM107\ & ( 
-- (\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM81\ & ((\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM85\) # (\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM83\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001110111000000000111011100010001111111110001000111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM83\,
	datab => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM85\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM81\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-2]_OTERM107\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-2]~13_combout\);

-- Location: LABCELL_X22_Y60_N45
\TheRxFsk|Bandpasses:4:Bandpass1|Add4~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add4~5_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass1|Sum\(0) ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed\(0) ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add4~66\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add4~6\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass1|Sum\(0) ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed\(0) ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add4~66\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111110000000000000000000000000101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum\(0),
	dataf => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed\(0),
	cin => \TheRxFsk|Bandpasses:4:Bandpass1|Add4~66\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass1|Add4~5_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass1|Add4~6\);

-- Location: FF_X19_Y59_N37
\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-3]_NEW_REG112\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~61_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-3]_OTERM113\);

-- Location: LABCELL_X19_Y60_N36
\TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-3]~12\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-3]~12_combout\ = (!\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM83\ & (\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM81\ & 
-- ((\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-3]_OTERM113\) # (\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM85\)))) # (\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM83\ & 
-- (((\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM85\ & \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-3]_OTERM113\)) # (\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM81\)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000101111111000000010111111100000001011111110000000101111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM83\,
	datab => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM85\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-3]_OTERM113\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM81\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-3]~12_combout\);

-- Location: FF_X19_Y59_N35
\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-4]_NEW_REG118\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~57_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-4]_OTERM119\);

-- Location: LABCELL_X19_Y60_N45
\TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-4]~11\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-4]~11_combout\ = (!\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM83\ & (\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM81\ & 
-- ((\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-4]_OTERM119\) # (\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM85\)))) # (\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM83\ & 
-- (((\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM85\ & \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-4]_OTERM119\)) # (\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM81\)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000101111111000000010111111100000001011111110000000101111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM83\,
	datab => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM85\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-4]_OTERM119\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM81\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-4]~11_combout\);

-- Location: FF_X19_Y59_N31
\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-5]_NEW_REG124\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~53_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-5]_OTERM125\);

-- Location: LABCELL_X19_Y60_N42
\TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-5]~10\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-5]~10_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-5]_OTERM125\ & ( ((\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM83\ & 
-- \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM85\)) # (\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM81\) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-5]_OTERM125\ & ( 
-- (\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM81\ & ((\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM85\) # (\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM83\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000011100000111000001110000011100011111000111110001111100011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM83\,
	datab => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM85\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM81\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-5]_OTERM125\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-5]~10_combout\);

-- Location: FF_X19_Y59_N28
\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-6]_NEW_REG130\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~49_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-6]_OTERM131\);

-- Location: LABCELL_X19_Y60_N27
\TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-6]~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-6]~9_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-6]_OTERM131\ & ( ((\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM83\ & 
-- \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM85\)) # (\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM81\) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-6]_OTERM131\ & ( 
-- (\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM81\ & ((\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM85\) # (\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM83\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001110111000000000111011100010001111111110001000111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM83\,
	datab => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM85\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM81\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-6]_OTERM131\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-6]~9_combout\);

-- Location: FF_X19_Y59_N26
\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-7]_NEW_REG136\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~45_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-7]_OTERM137\);

-- Location: LABCELL_X19_Y60_N24
\TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-7]~8\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-7]~8_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-7]_OTERM137\ & ( ((\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM83\ & 
-- \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM85\)) # (\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM81\) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-7]_OTERM137\ & ( 
-- (\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM81\ & ((\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM85\) # (\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM83\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000011100000111000001110000011100011111000111110001111100011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM83\,
	datab => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM85\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM81\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-7]_OTERM137\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-7]~8_combout\);

-- Location: FF_X19_Y59_N22
\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-8]_NEW_REG142\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~41_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-8]_OTERM143\);

-- Location: LABCELL_X19_Y60_N57
\TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-8]~7\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-8]~7_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-8]_OTERM143\ & ( ((\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM83\ & 
-- \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM85\)) # (\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM81\) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-8]_OTERM143\ & ( 
-- (\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM81\ & ((\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM85\) # (\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM83\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001110111000000000111011100010001111111110001000111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM83\,
	datab => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM85\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM81\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-8]_OTERM143\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-8]~7_combout\);

-- Location: FF_X19_Y59_N19
\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-9]_NEW_REG148\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~37_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-9]_OTERM149\);

-- Location: LABCELL_X19_Y60_N54
\TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-9]~6\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-9]~6_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-9]_OTERM149\ & ( ((\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM83\ & 
-- \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM85\)) # (\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM81\) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-9]_OTERM149\ & ( 
-- (\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM81\ & ((\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM85\) # (\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM83\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000011100000111000001110000011100011111000111110001111100011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM83\,
	datab => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM85\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM81\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-9]_OTERM149\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-9]~6_combout\);

-- Location: FF_X19_Y59_N16
\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-10]_NEW_REG154\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~33_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-10]_OTERM155\);

-- Location: LABCELL_X19_Y60_N15
\TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-10]~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-10]~5_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM83\ & ( \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-10]_OTERM155\ & ( 
-- (\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM85\) # (\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM81\) ) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM83\ & ( 
-- \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-10]_OTERM155\ & ( \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM81\ ) ) ) # ( \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM83\ & ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-10]_OTERM155\ & ( \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM81\ ) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM83\ & ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-10]_OTERM155\ & ( (\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM81\ & \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM85\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100000101010101010101010101010101010101010101111101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM81\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM85\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM83\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-10]_OTERM155\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-10]~5_combout\);

-- Location: FF_X19_Y59_N13
\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-11]_NEW_REG160\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~29_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-11]_OTERM161\);

-- Location: LABCELL_X19_Y60_N0
\TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-11]~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-11]~4_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-11]_OTERM161\ & ( ((\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM83\ & 
-- \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM85\)) # (\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM81\) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-11]_OTERM161\ & ( 
-- (\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM81\ & ((\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM85\) # (\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM83\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000011100000111000001110000011100011111000111110001111100011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM83\,
	datab => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM85\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM81\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-11]_OTERM161\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-11]~4_combout\);

-- Location: FF_X19_Y59_N10
\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-12]_NEW_REG166\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~25_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-12]_OTERM167\);

-- Location: LABCELL_X19_Y60_N9
\TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-12]~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-12]~3_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM83\ & ( ((\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM85\ & 
-- \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-12]_OTERM167\)) # (\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM81\) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM83\ & ( 
-- (\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM81\ & ((\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-12]_OTERM167\) # (\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM85\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010101010101010101010101111100000101010101010101010101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM81\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM85\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-12]_OTERM167\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM83\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-12]~3_combout\);

-- Location: FF_X19_Y59_N7
\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-13]_NEW_REG172\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~21_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-13]_OTERM173\);

-- Location: LABCELL_X19_Y60_N48
\TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-13]~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-13]~2_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM83\ & ( \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-13]_OTERM173\ & ( 
-- (\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM81\) # (\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM85\) ) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM83\ & ( 
-- \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-13]_OTERM173\ & ( \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM81\ ) ) ) # ( \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM83\ & ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-13]_OTERM173\ & ( \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM81\ ) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM83\ & ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-13]_OTERM173\ & ( (\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM85\ & \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM81\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100000011000011110000111100001111000011110011111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM85\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM81\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM83\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-13]_OTERM173\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-13]~2_combout\);

-- Location: FF_X19_Y59_N4
\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-14]_NEW_REG178\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~17_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-14]_OTERM179\);

-- Location: LABCELL_X19_Y60_N33
\TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-14]~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-14]~1_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM83\ & ( \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-14]_OTERM179\ & ( 
-- (\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM85\) # (\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM81\) ) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM83\ & ( 
-- \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-14]_OTERM179\ & ( \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM81\ ) ) ) # ( \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM83\ & ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-14]_OTERM179\ & ( \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM81\ ) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM83\ & ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-14]_OTERM179\ & ( (\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM81\ & \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM85\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100000101010101010101010101010101010101010101111101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM81\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM85\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM83\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-14]_OTERM179\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-14]~1_combout\);

-- Location: FF_X19_Y59_N2
\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_NEW_REG86\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass1|Add3~13_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM87\);

-- Location: LABCELL_X19_Y60_N3
\TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-15]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-15]~0_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM87\ & ( ((\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM83\ & 
-- \TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM85\)) # (\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM81\) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM87\ & ( 
-- (\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM81\ & ((\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM85\) # (\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed[-15]_OTERM83\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001110111000000000111011100010001111111110001000111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM83\,
	datab => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM85\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM81\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM87\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-15]~0_combout\);

-- Location: MLABCELL_X21_Y60_N42
\TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-15]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-15]~0_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-15]~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass1|Add4~5_sumout\ & ( (!\TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-15]~0_combout\) # 
-- (\TheRxFsk|Bandpasses:4:Bandpass1|Add4~1_sumout\) ) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass1|Sum[-15]~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass1|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-15]~0_combout\) # 
-- (\TheRxFsk|Bandpasses:4:Bandpass1|Add4~1_sumout\) ) ) ) # ( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-15]~q\ & ( !\TheRxFsk|Bandpasses:4:Bandpass1|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:4:Bandpass1|Add4~1_sumout\ & 
-- !\TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-15]~0_combout\) ) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass1|Sum[-15]~q\ & ( !\TheRxFsk|Bandpasses:4:Bandpass1|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:4:Bandpass1|Add4~1_sumout\ & 
-- \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-15]~0_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100000011001100000011000000111111001111111111001111110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~1_sumout\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResult[-15]~0_combout\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-15]~q\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~5_sumout\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-15]~0_combout\);

-- Location: FF_X16_Y62_N32
\TheRxFsk|Bandpasses:4:Bandpass1|R.SumState.SumValid\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	asdata => \TheRxFsk|Bandpasses:4:Bandpass1|R.SumState.SumWait2~q\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass1|R.SumState.SumValid~q\);

-- Location: LABCELL_X16_Y62_N42
\TheRxFsk|Bandpasses:4:Bandpass1|Selector0~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Selector0~0_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass1|R.SumState.Idle~q\ & ( \TheI2sToPar|ValL~q\ & ( !\TheRxFsk|Bandpasses:4:Bandpass1|R.SumState.SumValid~q\ ) ) ) # ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass1|R.SumState.Idle~q\ & ( \TheI2sToPar|ValL~q\ & ( !\TheRxFsk|Bandpasses:4:Bandpass1|R.SumState.SumValid~q\ ) ) ) # ( \TheRxFsk|Bandpasses:4:Bandpass1|R.SumState.Idle~q\ & ( !\TheI2sToPar|ValL~q\ & ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass1|R.SumState.SumValid~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111110000000011111111000000001111111100000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_R.SumState.SumValid~q\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_R.SumState.Idle~q\,
	dataf => \TheI2sToPar|ALT_INV_ValL~q\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|Selector0~0_combout\);

-- Location: FF_X16_Y62_N44
\TheRxFsk|Bandpasses:4:Bandpass1|R.SumState.Idle\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass1|Selector0~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass1|R.SumState.Idle~q\);

-- Location: LABCELL_X16_Y62_N27
\TheRxFsk|Bandpasses:4:Bandpass1|Selector1~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Selector1~0_combout\ = ( \TheI2sToPar|ValL~q\ & ( !\TheRxFsk|Bandpasses:4:Bandpass1|R.SumState.Idle~q\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011001100110011001100110011001100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_R.SumState.Idle~q\,
	dataf => \TheI2sToPar|ALT_INV_ValL~q\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|Selector1~0_combout\);

-- Location: FF_X16_Y62_N28
\TheRxFsk|Bandpasses:4:Bandpass1|R.SumState.SumEnable\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass1|Selector1~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass1|R.SumState.SumEnable~q\);

-- Location: LABCELL_X16_Y62_N12
\TheRxFsk|Bandpasses:4:Bandpass1|Selector2~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Selector2~0_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass1|R.SumState.SumEnable~q\ ) # ( !\TheRxFsk|Bandpasses:4:Bandpass1|R.SumState.SumEnable~q\ & ( (\TheRxFsk|Bandpasses:4:Bandpass1|R.SumState.SumSelect~q\ & 
-- ((!\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~1_combout\) # (!\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~0_combout\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011101110000000001110111011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:11:Bandpass1|ALT_INV_Equal1~1_combout\,
	datab => \TheRxFsk|Bandpasses:11:Bandpass1|ALT_INV_Equal1~0_combout\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_R.SumState.SumSelect~q\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_R.SumState.SumEnable~q\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|Selector2~0_combout\);

-- Location: FF_X16_Y62_N14
\TheRxFsk|Bandpasses:4:Bandpass1|R.SumState.SumSelect\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass1|Selector2~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass1|R.SumState.SumSelect~q\);

-- Location: LABCELL_X16_Y62_N15
\TheRxFsk|Bandpasses:4:Bandpass1|Selector3~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Selector3~0_combout\ = (\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~1_combout\ & (\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~0_combout\ & \TheRxFsk|Bandpasses:4:Bandpass1|R.SumState.SumSelect~q\))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000100000001000000010000000100000001000000010000000100000001",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:11:Bandpass1|ALT_INV_Equal1~1_combout\,
	datab => \TheRxFsk|Bandpasses:11:Bandpass1|ALT_INV_Equal1~0_combout\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_R.SumState.SumSelect~q\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|Selector3~0_combout\);

-- Location: FF_X16_Y62_N17
\TheRxFsk|Bandpasses:4:Bandpass1|R.SumState.SumWait1\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass1|Selector3~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass1|R.SumState.SumWait1~q\);

-- Location: FF_X16_Y62_N8
\TheRxFsk|Bandpasses:4:Bandpass1|R.SumState.SumWait2\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	asdata => \TheRxFsk|Bandpasses:4:Bandpass1|R.SumState.SumWait1~q\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass1|R.SumState.SumWait2~q\);

-- Location: LABCELL_X16_Y62_N57
\TheRxFsk|Bandpasses:4:Bandpass1|Selector6~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Selector6~0_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass1|R.SelSumUp~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass1|R.SumState.SumEnable~q\ ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass1|R.SelSumUp~q\ & ( 
-- \TheRxFsk|Bandpasses:4:Bandpass1|R.SumState.SumEnable~q\ ) ) # ( \TheRxFsk|Bandpasses:4:Bandpass1|R.SelSumUp~q\ & ( !\TheRxFsk|Bandpasses:4:Bandpass1|R.SumState.SumEnable~q\ & ( !\TheRxFsk|Bandpasses:4:Bandpass1|R.SumState.SumWait2~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000110011001100110011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_R.SumState.SumWait2~q\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_R.SelSumUp~q\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_R.SumState.SumEnable~q\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|Selector6~0_combout\);

-- Location: FF_X16_Y62_N58
\TheRxFsk|Bandpasses:4:Bandpass1|R.SelSumUp\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass1|Selector6~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass1|R.SelSumUp~q\);

-- Location: LABCELL_X16_Y62_N36
\TheRxFsk|Bandpasses:4:Bandpass1|Selector7~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Selector7~0_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass1|R.EnableSumUp~q\ & ( \TheI2sToPar|ValL~q\ & ( (!\TheRxFsk|Bandpasses:4:Bandpass1|R.SumState.Idle~q\) # (!\TheRxFsk|Bandpasses:4:Bandpass1|R.SumState.SumWait2~q\) ) 
-- ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass1|R.EnableSumUp~q\ & ( \TheI2sToPar|ValL~q\ & ( !\TheRxFsk|Bandpasses:4:Bandpass1|R.SumState.Idle~q\ ) ) ) # ( \TheRxFsk|Bandpasses:4:Bandpass1|R.EnableSumUp~q\ & ( !\TheI2sToPar|ValL~q\ & ( 
-- (!\TheRxFsk|Bandpasses:4:Bandpass1|R.SumState.Idle~q\) # (!\TheRxFsk|Bandpasses:4:Bandpass1|R.SumState.SumWait2~q\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111100110011001100110011001111111111001100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_R.SumState.Idle~q\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_R.SumState.SumWait2~q\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_R.EnableSumUp~q\,
	dataf => \TheI2sToPar|ALT_INV_ValL~q\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|Selector7~0_combout\);

-- Location: FF_X16_Y62_N37
\TheRxFsk|Bandpasses:4:Bandpass1|R.EnableSumUp\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass1|Selector7~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass1|R.EnableSumUp~q\);

-- Location: FF_X21_Y60_N43
\TheRxFsk|Bandpasses:4:Bandpass1|Sum[-15]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-15]~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:4:Bandpass1|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-15]~q\);

-- Location: LABCELL_X22_Y60_N0
\TheRxFsk|Bandpasses:4:Bandpass1|Add4~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add4~10\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-15]~0_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-15]~q\ ) + ( !VCC ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000110011001100110000000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-15]~q\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResult[-15]~0_combout\,
	cin => GND,
	cout => \TheRxFsk|Bandpasses:4:Bandpass1|Add4~10\);

-- Location: LABCELL_X22_Y60_N3
\TheRxFsk|Bandpasses:4:Bandpass1|Add4~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add4~13_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-14]~1_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-14]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add4~10\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add4~14\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-14]~1_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-14]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add4~10\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111110000000000000000000000000101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResult[-14]~1_combout\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-14]~q\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass1|Add4~10\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass1|Add4~13_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass1|Add4~14\);

-- Location: MLABCELL_X21_Y60_N51
\TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-14]~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-14]~1_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass1|Add4~1_sumout\ & ( \TheRxFsk|Bandpasses:4:Bandpass1|Add4~5_sumout\ ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass1|Add4~1_sumout\ & ( 
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add4~5_sumout\ & ( \TheRxFsk|Bandpasses:4:Bandpass1|Add4~13_sumout\ ) ) ) # ( \TheRxFsk|Bandpasses:4:Bandpass1|Add4~1_sumout\ & ( !\TheRxFsk|Bandpasses:4:Bandpass1|Add4~5_sumout\ & ( 
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add4~13_sumout\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000010101010101010101010101010101011111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~13_sumout\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~1_sumout\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~5_sumout\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-14]~1_combout\);

-- Location: FF_X21_Y60_N52
\TheRxFsk|Bandpasses:4:Bandpass1|Sum[-14]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-14]~1_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:4:Bandpass1|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-14]~q\);

-- Location: LABCELL_X22_Y60_N6
\TheRxFsk|Bandpasses:4:Bandpass1|Add4~17\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add4~17_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-13]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-13]~2_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add4~14\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add4~18\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-13]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-13]~2_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add4~14\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000110011001100110000000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResult[-13]~2_combout\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-13]~q\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass1|Add4~14\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass1|Add4~17_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass1|Add4~18\);

-- Location: MLABCELL_X21_Y60_N54
\TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-13]~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-13]~2_combout\ = (!\TheRxFsk|Bandpasses:4:Bandpass1|Add4~5_sumout\ & (\TheRxFsk|Bandpasses:4:Bandpass1|Add4~1_sumout\ & \TheRxFsk|Bandpasses:4:Bandpass1|Add4~17_sumout\)) # 
-- (\TheRxFsk|Bandpasses:4:Bandpass1|Add4~5_sumout\ & ((\TheRxFsk|Bandpasses:4:Bandpass1|Add4~17_sumout\) # (\TheRxFsk|Bandpasses:4:Bandpass1|Add4~1_sumout\)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001011100010111000101110001011100010111000101110001011100010111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~5_sumout\,
	datab => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~1_sumout\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~17_sumout\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-13]~2_combout\);

-- Location: FF_X21_Y60_N55
\TheRxFsk|Bandpasses:4:Bandpass1|Sum[-13]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-13]~2_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:4:Bandpass1|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-13]~q\);

-- Location: LABCELL_X22_Y60_N9
\TheRxFsk|Bandpasses:4:Bandpass1|Add4~21\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add4~21_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-12]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-12]~3_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add4~18\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add4~22\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-12]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-12]~3_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add4~18\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111110000000000000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-12]~q\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResult[-12]~3_combout\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass1|Add4~18\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass1|Add4~21_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass1|Add4~22\);

-- Location: MLABCELL_X21_Y60_N57
\TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-12]~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-12]~3_combout\ = (!\TheRxFsk|Bandpasses:4:Bandpass1|Add4~5_sumout\ & (\TheRxFsk|Bandpasses:4:Bandpass1|Add4~1_sumout\ & \TheRxFsk|Bandpasses:4:Bandpass1|Add4~21_sumout\)) # 
-- (\TheRxFsk|Bandpasses:4:Bandpass1|Add4~5_sumout\ & ((\TheRxFsk|Bandpasses:4:Bandpass1|Add4~21_sumout\) # (\TheRxFsk|Bandpasses:4:Bandpass1|Add4~1_sumout\)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000101110111000100010111011100010001011101110001000101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~5_sumout\,
	datab => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~1_sumout\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~21_sumout\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-12]~3_combout\);

-- Location: FF_X21_Y60_N58
\TheRxFsk|Bandpasses:4:Bandpass1|Sum[-12]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-12]~3_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:4:Bandpass1|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-12]~q\);

-- Location: LABCELL_X22_Y60_N12
\TheRxFsk|Bandpasses:4:Bandpass1|Add4~25\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add4~25_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-11]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-11]~4_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add4~22\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add4~26\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-11]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-11]~4_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add4~22\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResult[-11]~4_combout\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-11]~q\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass1|Add4~22\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass1|Add4~25_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass1|Add4~26\);

-- Location: MLABCELL_X21_Y60_N12
\TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-11]~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-11]~4_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass1|Add4~25_sumout\ & ( (\TheRxFsk|Bandpasses:4:Bandpass1|Add4~1_sumout\) # (\TheRxFsk|Bandpasses:4:Bandpass1|Add4~5_sumout\) ) ) # ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass1|Add4~25_sumout\ & ( (\TheRxFsk|Bandpasses:4:Bandpass1|Add4~5_sumout\ & \TheRxFsk|Bandpasses:4:Bandpass1|Add4~1_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000100010001000100010001000101110111011101110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~5_sumout\,
	datab => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~1_sumout\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~25_sumout\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-11]~4_combout\);

-- Location: FF_X21_Y60_N13
\TheRxFsk|Bandpasses:4:Bandpass1|Sum[-11]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-11]~4_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:4:Bandpass1|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-11]~q\);

-- Location: LABCELL_X22_Y60_N15
\TheRxFsk|Bandpasses:4:Bandpass1|Add4~29\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add4~29_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-10]~5_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-10]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add4~26\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add4~30\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-10]~5_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-10]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add4~26\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111110000000000000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResult[-10]~5_combout\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-10]~q\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass1|Add4~26\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass1|Add4~29_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass1|Add4~30\);

-- Location: MLABCELL_X21_Y60_N15
\TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-10]~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-10]~5_combout\ = (!\TheRxFsk|Bandpasses:4:Bandpass1|Add4~5_sumout\ & (\TheRxFsk|Bandpasses:4:Bandpass1|Add4~1_sumout\ & \TheRxFsk|Bandpasses:4:Bandpass1|Add4~29_sumout\)) # 
-- (\TheRxFsk|Bandpasses:4:Bandpass1|Add4~5_sumout\ & ((\TheRxFsk|Bandpasses:4:Bandpass1|Add4~29_sumout\) # (\TheRxFsk|Bandpasses:4:Bandpass1|Add4~1_sumout\)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000101110111000100010111011100010001011101110001000101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~5_sumout\,
	datab => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~1_sumout\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~29_sumout\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-10]~5_combout\);

-- Location: FF_X21_Y60_N16
\TheRxFsk|Bandpasses:4:Bandpass1|Sum[-10]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-10]~5_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:4:Bandpass1|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-10]~q\);

-- Location: LABCELL_X22_Y60_N18
\TheRxFsk|Bandpasses:4:Bandpass1|Add4~33\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add4~33_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-9]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-9]~6_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add4~30\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add4~34\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-9]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-9]~6_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add4~30\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000101010101010101000000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResult[-9]~6_combout\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-9]~q\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass1|Add4~30\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass1|Add4~33_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass1|Add4~34\);

-- Location: MLABCELL_X21_Y60_N18
\TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-9]~6\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-9]~6_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass1|Add4~33_sumout\ & ( (\TheRxFsk|Bandpasses:4:Bandpass1|Add4~1_sumout\) # (\TheRxFsk|Bandpasses:4:Bandpass1|Add4~5_sumout\) ) ) # ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass1|Add4~33_sumout\ & ( (\TheRxFsk|Bandpasses:4:Bandpass1|Add4~5_sumout\ & \TheRxFsk|Bandpasses:4:Bandpass1|Add4~1_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000100010001000100010001000101110111011101110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~5_sumout\,
	datab => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~1_sumout\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~33_sumout\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-9]~6_combout\);

-- Location: FF_X21_Y60_N19
\TheRxFsk|Bandpasses:4:Bandpass1|Sum[-9]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-9]~6_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:4:Bandpass1|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-9]~q\);

-- Location: LABCELL_X22_Y60_N21
\TheRxFsk|Bandpasses:4:Bandpass1|Add4~37\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add4~37_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-8]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-8]~7_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add4~34\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add4~38\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-8]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-8]~7_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add4~34\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResult[-8]~7_combout\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-8]~q\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass1|Add4~34\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass1|Add4~37_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass1|Add4~38\);

-- Location: MLABCELL_X21_Y60_N21
\TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-8]~7\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-8]~7_combout\ = (!\TheRxFsk|Bandpasses:4:Bandpass1|Add4~5_sumout\ & (\TheRxFsk|Bandpasses:4:Bandpass1|Add4~1_sumout\ & \TheRxFsk|Bandpasses:4:Bandpass1|Add4~37_sumout\)) # 
-- (\TheRxFsk|Bandpasses:4:Bandpass1|Add4~5_sumout\ & ((\TheRxFsk|Bandpasses:4:Bandpass1|Add4~37_sumout\) # (\TheRxFsk|Bandpasses:4:Bandpass1|Add4~1_sumout\)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000101110111000100010111011100010001011101110001000101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~5_sumout\,
	datab => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~1_sumout\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~37_sumout\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-8]~7_combout\);

-- Location: FF_X21_Y60_N22
\TheRxFsk|Bandpasses:4:Bandpass1|Sum[-8]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-8]~7_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:4:Bandpass1|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-8]~q\);

-- Location: LABCELL_X22_Y60_N24
\TheRxFsk|Bandpasses:4:Bandpass1|Add4~41\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add4~41_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-7]~8_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-7]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add4~38\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add4~42\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-7]~8_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-7]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add4~38\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111110000000000000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResult[-7]~8_combout\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-7]~q\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass1|Add4~38\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass1|Add4~41_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass1|Add4~42\);

-- Location: MLABCELL_X21_Y60_N24
\TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-7]~8\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-7]~8_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass1|Add4~41_sumout\ & ( (\TheRxFsk|Bandpasses:4:Bandpass1|Add4~1_sumout\) # (\TheRxFsk|Bandpasses:4:Bandpass1|Add4~5_sumout\) ) ) # ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass1|Add4~41_sumout\ & ( (\TheRxFsk|Bandpasses:4:Bandpass1|Add4~5_sumout\ & \TheRxFsk|Bandpasses:4:Bandpass1|Add4~1_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000100010001000100010001000101110111011101110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~5_sumout\,
	datab => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~1_sumout\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~41_sumout\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-7]~8_combout\);

-- Location: FF_X21_Y60_N25
\TheRxFsk|Bandpasses:4:Bandpass1|Sum[-7]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-7]~8_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:4:Bandpass1|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-7]~q\);

-- Location: LABCELL_X22_Y60_N27
\TheRxFsk|Bandpasses:4:Bandpass1|Add4~45\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add4~45_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-6]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-6]~9_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add4~42\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add4~46\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-6]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-6]~9_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add4~42\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-6]~q\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResult[-6]~9_combout\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass1|Add4~42\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass1|Add4~45_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass1|Add4~46\);

-- Location: MLABCELL_X21_Y60_N27
\TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-6]~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-6]~9_combout\ = (!\TheRxFsk|Bandpasses:4:Bandpass1|Add4~5_sumout\ & (\TheRxFsk|Bandpasses:4:Bandpass1|Add4~1_sumout\ & \TheRxFsk|Bandpasses:4:Bandpass1|Add4~45_sumout\)) # 
-- (\TheRxFsk|Bandpasses:4:Bandpass1|Add4~5_sumout\ & ((\TheRxFsk|Bandpasses:4:Bandpass1|Add4~45_sumout\) # (\TheRxFsk|Bandpasses:4:Bandpass1|Add4~1_sumout\)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000101110111000100010111011100010001011101110001000101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~5_sumout\,
	datab => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~1_sumout\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~45_sumout\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-6]~9_combout\);

-- Location: FF_X21_Y60_N28
\TheRxFsk|Bandpasses:4:Bandpass1|Sum[-6]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-6]~9_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:4:Bandpass1|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-6]~q\);

-- Location: LABCELL_X22_Y60_N30
\TheRxFsk|Bandpasses:4:Bandpass1|Add4~49\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add4~49_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-5]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-5]~10_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add4~46\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add4~50\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-5]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-5]~10_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add4~46\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000110011001100110000000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResult[-5]~10_combout\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-5]~q\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass1|Add4~46\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass1|Add4~49_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass1|Add4~50\);

-- Location: MLABCELL_X21_Y60_N30
\TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-5]~10\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-5]~10_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass1|Add4~49_sumout\ & ( (\TheRxFsk|Bandpasses:4:Bandpass1|Add4~1_sumout\) # (\TheRxFsk|Bandpasses:4:Bandpass1|Add4~5_sumout\) ) ) # ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass1|Add4~49_sumout\ & ( (\TheRxFsk|Bandpasses:4:Bandpass1|Add4~5_sumout\ & \TheRxFsk|Bandpasses:4:Bandpass1|Add4~1_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000100010001000100010001000101110111011101110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~5_sumout\,
	datab => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~1_sumout\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~49_sumout\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-5]~10_combout\);

-- Location: FF_X21_Y60_N31
\TheRxFsk|Bandpasses:4:Bandpass1|Sum[-5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-5]~10_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:4:Bandpass1|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-5]~q\);

-- Location: LABCELL_X22_Y60_N33
\TheRxFsk|Bandpasses:4:Bandpass1|Add4~53\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add4~53_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-4]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-4]~11_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add4~50\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add4~54\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-4]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-4]~11_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add4~50\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-4]~q\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResult[-4]~11_combout\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass1|Add4~50\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass1|Add4~53_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass1|Add4~54\);

-- Location: MLABCELL_X21_Y60_N33
\TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-4]~11\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-4]~11_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass1|Add4~53_sumout\ & ( (\TheRxFsk|Bandpasses:4:Bandpass1|Add4~1_sumout\) # (\TheRxFsk|Bandpasses:4:Bandpass1|Add4~5_sumout\) ) ) # ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass1|Add4~53_sumout\ & ( (\TheRxFsk|Bandpasses:4:Bandpass1|Add4~5_sumout\ & \TheRxFsk|Bandpasses:4:Bandpass1|Add4~1_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000100010001000100010001000101110111011101110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~5_sumout\,
	datab => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~1_sumout\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~53_sumout\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-4]~11_combout\);

-- Location: FF_X21_Y60_N34
\TheRxFsk|Bandpasses:4:Bandpass1|Sum[-4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-4]~11_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:4:Bandpass1|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-4]~q\);

-- Location: LABCELL_X22_Y60_N36
\TheRxFsk|Bandpasses:4:Bandpass1|Add4~57\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add4~57_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-3]~12_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-3]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add4~54\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add4~58\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-3]~12_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-3]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add4~54\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111110000000000000000000000000011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResult[-3]~12_combout\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-3]~q\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass1|Add4~54\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass1|Add4~57_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass1|Add4~58\);

-- Location: MLABCELL_X21_Y60_N0
\TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-3]~12\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-3]~12_combout\ = (!\TheRxFsk|Bandpasses:4:Bandpass1|Add4~5_sumout\ & (\TheRxFsk|Bandpasses:4:Bandpass1|Add4~1_sumout\ & \TheRxFsk|Bandpasses:4:Bandpass1|Add4~57_sumout\)) # 
-- (\TheRxFsk|Bandpasses:4:Bandpass1|Add4~5_sumout\ & ((\TheRxFsk|Bandpasses:4:Bandpass1|Add4~57_sumout\) # (\TheRxFsk|Bandpasses:4:Bandpass1|Add4~1_sumout\)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000101110111000100010111011100010001011101110001000101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~5_sumout\,
	datab => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~1_sumout\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~57_sumout\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-3]~12_combout\);

-- Location: FF_X21_Y60_N1
\TheRxFsk|Bandpasses:4:Bandpass1|Sum[-3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-3]~12_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:4:Bandpass1|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-3]~q\);

-- Location: LABCELL_X22_Y60_N39
\TheRxFsk|Bandpasses:4:Bandpass1|Add4~61\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add4~61_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-2]~13_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-2]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add4~58\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add4~62\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-2]~13_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-2]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add4~58\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111110000000000000000000000000101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResult[-2]~13_combout\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-2]~q\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass1|Add4~58\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass1|Add4~61_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass1|Add4~62\);

-- Location: MLABCELL_X21_Y60_N3
\TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-2]~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-2]~13_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass1|Add4~61_sumout\ & ( (\TheRxFsk|Bandpasses:4:Bandpass1|Add4~1_sumout\) # (\TheRxFsk|Bandpasses:4:Bandpass1|Add4~5_sumout\) ) ) # ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass1|Add4~61_sumout\ & ( (\TheRxFsk|Bandpasses:4:Bandpass1|Add4~5_sumout\ & \TheRxFsk|Bandpasses:4:Bandpass1|Add4~1_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000100010001000100010001000101110111011101110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~5_sumout\,
	datab => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~1_sumout\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~61_sumout\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-2]~13_combout\);

-- Location: FF_X21_Y60_N4
\TheRxFsk|Bandpasses:4:Bandpass1|Sum[-2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-2]~13_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:4:Bandpass1|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-2]~q\);

-- Location: LABCELL_X22_Y60_N42
\TheRxFsk|Bandpasses:4:Bandpass1|Add4~65\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add4~65_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-1]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-1]~14_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add4~62\ ))
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add4~66\ = CARRY(( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-1]~q\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|MultResult[-1]~14_combout\ ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add4~62\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000110011001100110000000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResult[-1]~14_combout\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-1]~q\,
	cin => \TheRxFsk|Bandpasses:4:Bandpass1|Add4~62\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass1|Add4~65_sumout\,
	cout => \TheRxFsk|Bandpasses:4:Bandpass1|Add4~66\);

-- Location: MLABCELL_X21_Y60_N9
\TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-1]~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-1]~14_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass1|Add4~1_sumout\ & ( \TheRxFsk|Bandpasses:4:Bandpass1|Add4~5_sumout\ ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass1|Add4~1_sumout\ & ( 
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add4~5_sumout\ & ( \TheRxFsk|Bandpasses:4:Bandpass1|Add4~65_sumout\ ) ) ) # ( \TheRxFsk|Bandpasses:4:Bandpass1|Add4~1_sumout\ & ( !\TheRxFsk|Bandpasses:4:Bandpass1|Add4~5_sumout\ & ( 
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add4~65_sumout\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000011110000111100001111000011111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~65_sumout\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~1_sumout\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~5_sumout\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-1]~14_combout\);

-- Location: FF_X21_Y60_N10
\TheRxFsk|Bandpasses:4:Bandpass1|Sum[-1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass1|NextSum[-1]~14_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:4:Bandpass1|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-1]~q\);

-- Location: LABCELL_X22_Y60_N48
\TheRxFsk|Bandpasses:4:Bandpass1|Add4~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add4~1_sumout\ = SUM(( \TheRxFsk|Bandpasses:4:Bandpass1|Sum\(0) ) + ( !\TheRxFsk|Bandpasses:4:Bandpass1|MultResultDelayed\(0) ) + ( \TheRxFsk|Bandpasses:4:Bandpass1|Add4~6\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000010101010101010100000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_MultResultDelayed\(0),
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum\(0),
	cin => \TheRxFsk|Bandpasses:4:Bandpass1|Add4~6\,
	sumout => \TheRxFsk|Bandpasses:4:Bandpass1|Add4~1_sumout\);

-- Location: MLABCELL_X21_Y60_N36
\TheRxFsk|Bandpasses:4:Bandpass1|Add4~1_wirecell\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:4:Bandpass1|Add4~1_wirecell_combout\ = ( !\TheRxFsk|Bandpasses:4:Bandpass1|Add4~1_sumout\ )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111111111111000000000000000011111111111111110000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datae => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Add4~1_sumout\,
	combout => \TheRxFsk|Bandpasses:4:Bandpass1|Add4~1_wirecell_combout\);

-- Location: FF_X21_Y60_N37
\TheRxFsk|Bandpasses:4:Bandpass1|Sum[0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:4:Bandpass1|Add4~1_wirecell_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:4:Bandpass1|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass1|Sum\(0));

-- Location: MLABCELL_X15_Y61_N42
\TheRxFsk|Bandpasses:7:Bandpass1|Sample[-15]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-15]~0_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a0\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-15]~q\) # (\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\) ) 
-- ) # ( !\TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a0\ & ( (!\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-15]~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011110000000000001111000000001111111111110000111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-15]~q\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a0\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-15]~0_combout\);

-- Location: LABCELL_X17_Y61_N36
\TheRxFsk|Bandpasses:7:Bandpass1|Sample[-14]~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-14]~1_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a1\ ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & 
-- ( \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a1\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-14]~q\ ) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( 
-- !\TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a1\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-14]~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111000000000000000000001111000011111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-14]~q\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a1\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-14]~1_combout\);

-- Location: LABCELL_X17_Y61_N33
\TheRxFsk|Bandpasses:7:Bandpass1|Sample[-13]~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-13]~2_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a2\ ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & 
-- ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-13]~q\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010101010101000000001111111101010101010101010000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-13]~q\,
	datad => \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a2\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-13]~2_combout\);

-- Location: LABCELL_X17_Y63_N51
\TheRxFsk|Bandpasses:7:Bandpass1|Sample[-12]~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-12]~3_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a3\ ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & 
-- ( \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a3\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-12]~q\ ) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( 
-- !\TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a3\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-12]~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111000000000000000000001111000011111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-12]~q\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a3\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-12]~3_combout\);

-- Location: LABCELL_X17_Y63_N45
\TheRxFsk|Bandpasses:7:Bandpass1|Sample[-11]~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-11]~4_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-11]~q\ & ( \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a4\ ) ) # ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-11]~q\ & ( \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a4\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ ) ) ) # ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-11]~q\ 
-- & ( !\TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a4\ & ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000101010101010101001010101010101011111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-11]~q\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a4\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-11]~4_combout\);

-- Location: LABCELL_X16_Y63_N39
\TheRxFsk|Bandpasses:7:Bandpass1|Sample[-10]~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-10]~5_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a5\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\) # (\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-10]~q\) ) 
-- ) # ( !\TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a5\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-10]~q\ & !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100000000000011110000000000001111111111110000111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-10]~q\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a5\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-10]~5_combout\);

-- Location: LABCELL_X19_Y63_N39
\TheRxFsk|Bandpasses:7:Bandpass1|Sample[-9]~6\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-9]~6_combout\ = (!\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ((\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-9]~q\))) # (\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & 
-- (\TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a6\))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010110101111000001011010111100000101101011110000010110101111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a6\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-9]~q\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-9]~6_combout\);

-- Location: LABCELL_X18_Y62_N27
\TheRxFsk|Bandpasses:7:Bandpass1|Sample[-8]~7\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-8]~7_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a7\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\) # (\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-8]~q\) ) ) 
-- # ( !\TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a7\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-8]~q\ & !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101000001010000010100000101000001011111010111110101111101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-8]~q\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a7\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-8]~7_combout\);

-- Location: LABCELL_X16_Y63_N21
\TheRxFsk|Bandpasses:7:Bandpass1|Sample[-7]~8\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-7]~8_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a8\ ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & 
-- ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-7]~q\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010101010101000011110000111101010101010101010000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-7]~q\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a8\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-7]~8_combout\);

-- Location: MLABCELL_X15_Y63_N33
\TheRxFsk|Bandpasses:7:Bandpass1|Sample[-6]~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-6]~9_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-6]~q\ & ( (!\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\) # (\TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a9\) ) 
-- ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-6]~q\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a9\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001010101101010101111111100000000010101011010101011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	datad => \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a9\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-6]~q\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-6]~9_combout\);

-- Location: LABCELL_X16_Y61_N18
\TheRxFsk|Bandpasses:7:Bandpass1|Sample[-5]~10\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-5]~10_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-5]~q\ & ( \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a10\ ) ) # ( 
-- !\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-5]~q\ & ( \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a10\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ ) ) ) # ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-5]~q\ 
-- & ( !\TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a10\ & ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000110011001100110000110011001100111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-5]~q\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a10\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-5]~10_combout\);

-- Location: LABCELL_X16_Y61_N51
\TheRxFsk|Bandpasses:7:Bandpass1|Sample[-4]~11\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-4]~11_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a11\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\) # (\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-4]~q\) ) 
-- ) # ( !\TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a11\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-4]~q\ & !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101000001010000010111110101111101010000010100000101111101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-4]~q\,
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	datae => \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a11\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-4]~11_combout\);

-- Location: MLABCELL_X15_Y63_N54
\TheRxFsk|Bandpasses:7:Bandpass1|Sample[-3]~12\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-3]~12_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-3]~q\ & ( \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a12\ ) ) 
-- ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-3]~q\ ) ) # ( \TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( !\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-3]~q\ & ( 
-- \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a12\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000011110000111111111111111111110000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a12\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-3]~q\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-3]~12_combout\);

-- Location: LABCELL_X16_Y63_N33
\TheRxFsk|Bandpasses:7:Bandpass1|Sample[-2]~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-2]~13_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-2]~q\ & ( (!\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\) # (\TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a13\) 
-- ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-2]~q\ & ( (\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a13\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100000101101011111010111100000101000001011010111110101111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a13\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-2]~q\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-2]~13_combout\);

-- Location: LABCELL_X17_Y63_N12
\TheRxFsk|Bandpasses:7:Bandpass1|Sample[-1]~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-1]~14_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a14\ ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ 
-- & ( \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a14\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-1]~q\ ) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( 
-- !\TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a14\ & ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[-1]~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111000000000000000000001111000011111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed[-1]~q\,
	datae => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a14\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|Sample[-1]~14_combout\);

-- Location: FF_X13_Y63_N38
\TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed[0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	asdata => \TheI2sToPar|D\(15),
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed\(0));

-- Location: LABCELL_X13_Y63_N0
\TheRxFsk|Bandpasses:7:Bandpass1|Sample[0]~15\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Sample[0]~15_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & ( \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ram_block1a15\ ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass0|R.FirstSample~q\ & 
-- ( \TheRxFsk|Bandpasses:4:Bandpass0|DdryDelayed\(0) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011111111000000001111111100001111000011110000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a15\,
	datad => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_DdryDelayed\(0),
	dataf => \TheRxFsk|Bandpasses:4:Bandpass0|ALT_INV_R.FirstSample~q\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|Sample[0]~15_combout\);

-- Location: DSP_X20_Y61_N0
\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8\ : cyclonev_mac
-- pragma translate_off
GENERIC MAP (
	accumulate_clock => "none",
	ax_clock => "none",
	ax_width => 18,
	ay_scan_in_clock => "none",
	ay_scan_in_width => 19,
	ay_use_scan_in => "false",
	az_clock => "none",
	bx_clock => "none",
	by_clock => "none",
	by_use_scan_in => "false",
	bz_clock => "none",
	coef_a_0 => 0,
	coef_a_1 => 0,
	coef_a_2 => 0,
	coef_a_3 => 0,
	coef_a_4 => 0,
	coef_a_5 => 0,
	coef_a_6 => 0,
	coef_a_7 => 0,
	coef_b_0 => 0,
	coef_b_1 => 0,
	coef_b_2 => 0,
	coef_b_3 => 0,
	coef_b_4 => 0,
	coef_b_5 => 0,
	coef_b_6 => 0,
	coef_b_7 => 0,
	coef_sel_a_clock => "none",
	coef_sel_b_clock => "none",
	delay_scan_out_ay => "false",
	delay_scan_out_by => "false",
	enable_double_accum => "false",
	load_const_clock => "none",
	load_const_value => 0,
	mode_sub_location => 0,
	negate_clock => "none",
	operand_source_max => "input",
	operand_source_may => "input",
	operand_source_mbx => "input",
	operand_source_mby => "input",
	operation_mode => "m18x18_full",
	output_clock => "none",
	preadder_subtract_a => "false",
	preadder_subtract_b => "false",
	result_a_width => 64,
	signed_max => "true",
	signed_may => "true",
	signed_mbx => "false",
	signed_mby => "false",
	sub_clock => "none",
	use_chainadder => "false")
-- pragma translate_on
PORT MAP (
	sub => GND,
	negate => GND,
	ax => \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_AX_bus\,
	ay => \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_AY_bus\,
	resulta => \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_RESULTA_bus\);

-- Location: LABCELL_X19_Y61_N54
\TheRxFsk|Bandpasses:7:Bandpass1|vAdd~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|vAdd~1_combout\ = ( !\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~14\ & ( !\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~9\ & ( (!\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~15\ & (!\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~18\ & 
-- (!\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~17\ & !\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~16\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1000000000000000000000000000000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~15\,
	datab => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~18\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~17\,
	datad => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~16\,
	datae => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~14\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~9\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|vAdd~1_combout\);

-- Location: LABCELL_X18_Y61_N15
\TheRxFsk|Bandpasses:7:Bandpass1|vAdd~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|vAdd~2_combout\ = ( !\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~10\ & ( !\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~8_resulta\ & ( (!\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~11\ & (!\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~12\ & 
-- !\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~21\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1010000000000000000000000000000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~11\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~12\,
	datad => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~21\,
	datae => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~10\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~8_resulta\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|vAdd~2_combout\);

-- Location: LABCELL_X18_Y61_N27
\TheRxFsk|Bandpasses:7:Bandpass1|vAdd~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|vAdd~0_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~13\ & ( \TheRxFsk|Bandpasses:7:Bandpass1|vAdd~2_combout\ ) ) # ( !\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~13\ & ( \TheRxFsk|Bandpasses:7:Bandpass1|vAdd~2_combout\ & 
-- ( ((!\TheRxFsk|Bandpasses:7:Bandpass1|vAdd~1_combout\) # ((\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~20\) # (\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~22\))) # (\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~19\) ) ) ) # ( \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~13\ & ( 
-- !\TheRxFsk|Bandpasses:7:Bandpass1|vAdd~2_combout\ ) ) # ( !\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~13\ & ( !\TheRxFsk|Bandpasses:7:Bandpass1|vAdd~2_combout\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111111111111111111111111111111011111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~19\,
	datab => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_vAdd~1_combout\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~22\,
	datad => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~20\,
	datae => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~13\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_vAdd~2_combout\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|vAdd~0_combout\);

-- Location: LABCELL_X19_Y61_N0
\TheRxFsk|Bandpasses:7:Bandpass1|Add3~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add3~13_sumout\ = SUM(( (\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~39\ & \TheRxFsk|Bandpasses:7:Bandpass1|vAdd~0_combout\) ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~23\ ) + ( !VCC ))
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add3~14\ = CARRY(( (\TheRxFsk|Bandpasses:7:Bandpass1|Mult0~39\ & \TheRxFsk|Bandpasses:7:Bandpass1|vAdd~0_combout\) ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~23\ ) + ( !VCC ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~39\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~23\,
	datad => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_vAdd~0_combout\,
	cin => GND,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~13_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~14\);

-- Location: LABCELL_X19_Y61_N3
\TheRxFsk|Bandpasses:7:Bandpass1|Add3~17\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add3~17_sumout\ = SUM(( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~24\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add3~14\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add3~18\ = CARRY(( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~24\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add3~14\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~24\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~14\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~17_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~18\);

-- Location: LABCELL_X19_Y61_N6
\TheRxFsk|Bandpasses:7:Bandpass1|Add3~21\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add3~21_sumout\ = SUM(( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~25\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add3~18\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add3~22\ = CARRY(( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~25\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add3~18\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~25\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~18\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~21_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~22\);

-- Location: LABCELL_X19_Y61_N9
\TheRxFsk|Bandpasses:7:Bandpass1|Add3~25\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add3~25_sumout\ = SUM(( \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~26\ ) + ( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add3~22\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add3~26\ = CARRY(( \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~26\ ) + ( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add3~22\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~26\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~22\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~25_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~26\);

-- Location: LABCELL_X19_Y61_N12
\TheRxFsk|Bandpasses:7:Bandpass1|Add3~29\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add3~29_sumout\ = SUM(( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~27\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add3~26\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add3~30\ = CARRY(( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~27\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add3~26\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~27\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~26\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~29_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~30\);

-- Location: LABCELL_X19_Y61_N15
\TheRxFsk|Bandpasses:7:Bandpass1|Add3~33\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add3~33_sumout\ = SUM(( \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~28\ ) + ( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add3~30\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add3~34\ = CARRY(( \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~28\ ) + ( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add3~30\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~28\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~30\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~33_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~34\);

-- Location: LABCELL_X19_Y61_N18
\TheRxFsk|Bandpasses:7:Bandpass1|Add3~37\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add3~37_sumout\ = SUM(( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~29\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add3~34\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add3~38\ = CARRY(( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~29\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add3~34\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~29\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~34\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~37_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~38\);

-- Location: LABCELL_X19_Y61_N21
\TheRxFsk|Bandpasses:7:Bandpass1|Add3~41\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add3~41_sumout\ = SUM(( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~30\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add3~38\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add3~42\ = CARRY(( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~30\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add3~38\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~30\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~38\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~41_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~42\);

-- Location: LABCELL_X19_Y61_N24
\TheRxFsk|Bandpasses:7:Bandpass1|Add3~45\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add3~45_sumout\ = SUM(( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~31\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add3~42\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add3~46\ = CARRY(( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~31\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add3~42\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~31\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~42\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~45_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~46\);

-- Location: LABCELL_X19_Y61_N27
\TheRxFsk|Bandpasses:7:Bandpass1|Add3~49\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add3~49_sumout\ = SUM(( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~32\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add3~46\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add3~50\ = CARRY(( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~32\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add3~46\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~32\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~46\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~49_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~50\);

-- Location: LABCELL_X19_Y61_N30
\TheRxFsk|Bandpasses:7:Bandpass1|Add3~53\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add3~53_sumout\ = SUM(( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~33\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add3~50\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add3~54\ = CARRY(( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~33\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add3~50\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~33\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~50\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~53_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~54\);

-- Location: LABCELL_X19_Y61_N33
\TheRxFsk|Bandpasses:7:Bandpass1|Add3~57\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add3~57_sumout\ = SUM(( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~34\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add3~54\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add3~58\ = CARRY(( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~34\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add3~54\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~34\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~54\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~57_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~58\);

-- Location: LABCELL_X19_Y61_N36
\TheRxFsk|Bandpasses:7:Bandpass1|Add3~61\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add3~61_sumout\ = SUM(( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~35\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add3~58\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add3~62\ = CARRY(( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~35\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add3~58\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~35\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~58\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~61_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~62\);

-- Location: LABCELL_X19_Y61_N39
\TheRxFsk|Bandpasses:7:Bandpass1|Add3~65\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add3~65_sumout\ = SUM(( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~36\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add3~62\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add3~66\ = CARRY(( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~36\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add3~62\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000101010101010101000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~36\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~62\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~65_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~66\);

-- Location: LABCELL_X19_Y61_N42
\TheRxFsk|Bandpasses:7:Bandpass1|Add3~69\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add3~69_sumout\ = SUM(( \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~37\ ) + ( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add3~66\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add3~70\ = CARRY(( \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~37\ ) + ( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add3~66\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~37\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~66\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~69_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~70\);

-- Location: LABCELL_X19_Y61_N45
\TheRxFsk|Bandpasses:7:Bandpass1|Add3~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add3~9_sumout\ = SUM(( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~38\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add3~70\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add3~10\ = CARRY(( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~38\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add3~70\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000101010101010101000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~38\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~70\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~9_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~10\);

-- Location: LABCELL_X19_Y61_N48
\TheRxFsk|Bandpasses:7:Bandpass1|Add3~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add3~5_sumout\ = SUM(( \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~39\ ) + ( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add3~10\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add3~6\ = CARRY(( \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~39\ ) + ( GND ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add3~10\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~39\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~10\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~5_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~6\);

-- Location: LABCELL_X19_Y61_N51
\TheRxFsk|Bandpasses:7:Bandpass1|Add3~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add3~1_sumout\ = SUM(( VCC ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Mult0~39\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add3~6\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000001111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Mult0~39\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~6\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~1_sumout\);

-- Location: MLABCELL_X15_Y61_N30
\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[0]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[0]~0_combout\ = ( !\TheRxFsk|Bandpasses:7:Bandpass1|Add3~1_sumout\ )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111111111111111111111111111100000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add3~1_sumout\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[0]~0_combout\);

-- Location: FF_X15_Y61_N31
\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[0]~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed\(0));

-- Location: FF_X19_Y61_N47
\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_NEW_REG12\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~9_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM13\);

-- Location: FF_X19_Y61_N49
\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_NEW_REG10\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~5_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM11\);

-- Location: FF_X19_Y61_N53
\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_NEW_REG8\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~1_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM9\);

-- Location: FF_X19_Y61_N44
\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-1]_NEW_REG16\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~69_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-1]_OTERM17\);

-- Location: MLABCELL_X15_Y61_N21
\TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-1]~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-1]~14_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-1]_OTERM17\ & ( ((\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM13\ & 
-- \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM11\)) # (\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM9\) ) ) # ( !\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-1]_OTERM17\ & ( 
-- (\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM9\ & ((\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM11\) # (\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM13\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000011100000111000001110000011100011111000111110001111100011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM13\,
	datab => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM11\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM9\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-1]_OTERM17\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-1]~14_combout\);

-- Location: LABCELL_X17_Y62_N45
\TheRxFsk|Bandpasses:7:Bandpass1|Add4~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add4~5_sumout\ = SUM(( \TheRxFsk|Bandpasses:7:Bandpass1|Sum\(0) ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed\(0) ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add4~66\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add4~6\ = CARRY(( \TheRxFsk|Bandpasses:7:Bandpass1|Sum\(0) ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed\(0) ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add4~66\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111110000000000000000000000000101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum\(0),
	dataf => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed\(0),
	cin => \TheRxFsk|Bandpasses:7:Bandpass1|Add4~66\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass1|Add4~5_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass1|Add4~6\);

-- Location: FF_X19_Y61_N40
\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-2]_NEW_REG20\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~65_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-2]_OTERM21\);

-- Location: MLABCELL_X15_Y61_N48
\TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-2]~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-2]~13_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM13\ & ( ((\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM11\ & 
-- \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-2]_OTERM21\)) # (\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM9\) ) ) # ( !\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM13\ & ( 
-- (\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM9\ & ((\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-2]_OTERM21\) # (\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM11\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001011111000000000101111100000101111111110000010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM11\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-2]_OTERM21\,
	datad => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM9\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM13\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-2]~13_combout\);

-- Location: FF_X19_Y61_N37
\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-3]_NEW_REG24\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~61_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-3]_OTERM25\);

-- Location: MLABCELL_X15_Y61_N18
\TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-3]~12\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-3]~12_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-3]_OTERM25\ & ( ((\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM11\ & 
-- \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM13\)) # (\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM9\) ) ) # ( !\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-3]_OTERM25\ & ( 
-- (\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM9\ & ((\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM13\) # (\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM11\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000111111000000000011111100000011111111110000001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM11\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM13\,
	datad => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM9\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-3]_OTERM25\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-3]~12_combout\);

-- Location: FF_X19_Y61_N34
\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-4]_NEW_REG28\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~57_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-4]_OTERM29\);

-- Location: MLABCELL_X15_Y61_N27
\TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-4]~11\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-4]~11_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-4]_OTERM29\ & ( ((\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM13\ & 
-- \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM11\)) # (\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM9\) ) ) # ( !\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-4]_OTERM29\ & ( 
-- (\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM9\ & ((\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM11\) # (\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM13\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000011100000111000001110000011100011111000111110001111100011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM13\,
	datab => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM11\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM9\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-4]_OTERM29\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-4]~11_combout\);

-- Location: FF_X19_Y61_N32
\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-5]_NEW_REG32\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~53_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-5]_OTERM33\);

-- Location: MLABCELL_X15_Y61_N24
\TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-5]~10\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-5]~10_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-5]_OTERM33\ & ( ((\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM11\ & 
-- \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM13\)) # (\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM9\) ) ) # ( !\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-5]_OTERM33\ & ( 
-- (\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM9\ & ((\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM13\) # (\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM11\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000111111000000000011111100000011111111110000001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM11\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM13\,
	datad => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM9\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-5]_OTERM33\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-5]~10_combout\);

-- Location: FF_X19_Y61_N29
\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-6]_NEW_REG36\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~49_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-6]_OTERM37\);

-- Location: MLABCELL_X15_Y61_N57
\TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-6]~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-6]~9_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM13\ & ( ((\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM11\ & 
-- \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-6]_OTERM37\)) # (\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM9\) ) ) # ( !\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM13\ & ( 
-- (\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM9\ & ((\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-6]_OTERM37\) # (\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM11\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001001100010011000100110001001100110111001101110011011100110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM11\,
	datab => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM9\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-6]_OTERM37\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM13\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-6]~9_combout\);

-- Location: FF_X19_Y61_N25
\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-7]_NEW_REG42\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~45_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-7]_OTERM43\);

-- Location: MLABCELL_X15_Y61_N54
\TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-7]~8\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-7]~8_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM9\ & ( ((\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-7]_OTERM43\) # 
-- (\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM13\)) # (\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM11\) ) ) # ( !\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM9\ & ( 
-- (\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM11\ & (\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM13\ & \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-7]_OTERM43\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000101000000000000010101011111111111110101111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM11\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM13\,
	datad => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-7]_OTERM43\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM9\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-7]~8_combout\);

-- Location: FF_X19_Y61_N22
\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-8]_NEW_REG46\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~41_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-8]_OTERM47\);

-- Location: MLABCELL_X15_Y61_N45
\TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-8]~7\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-8]~7_combout\ = (!\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM13\ & (\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM9\ & 
-- ((\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-8]_OTERM47\) # (\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM11\)))) # (\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM13\ & 
-- (((\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM11\ & \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-8]_OTERM47\)) # (\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM9\)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000011100011111000001110001111100000111000111110000011100011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM13\,
	datab => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM11\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM9\,
	datad => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-8]_OTERM47\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-8]~7_combout\);

-- Location: FF_X19_Y61_N19
\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-9]_NEW_REG52\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~37_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-9]_OTERM53\);

-- Location: MLABCELL_X15_Y61_N51
\TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-9]~6\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-9]~6_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM13\ & ( ((\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM11\ & 
-- \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-9]_OTERM53\)) # (\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM9\) ) ) # ( !\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM13\ & ( 
-- (\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM9\ & ((\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-9]_OTERM53\) # (\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM11\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100001111000001010000111100001111010111110000111101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM11\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM9\,
	datad => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-9]_OTERM53\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM13\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-9]~6_combout\);

-- Location: FF_X19_Y61_N17
\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-10]_NEW_REG54\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~33_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-10]_OTERM55\);

-- Location: MLABCELL_X15_Y61_N3
\TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-10]~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-10]~5_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-10]_OTERM55\ & ( ((\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM13\ & 
-- \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM11\)) # (\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM9\) ) ) # ( !\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-10]_OTERM55\ & ( 
-- (\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM9\ & ((\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM11\) # (\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM13\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000011100000111000001110000011100011111000111110001111100011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM13\,
	datab => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM11\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM9\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-10]_OTERM55\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-10]~5_combout\);

-- Location: FF_X19_Y61_N13
\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-11]_NEW_REG58\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~29_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-11]_OTERM59\);

-- Location: MLABCELL_X15_Y61_N0
\TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-11]~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-11]~4_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-11]_OTERM59\ & ( ((\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM11\ & 
-- \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM13\)) # (\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM9\) ) ) # ( !\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-11]_OTERM59\ & ( 
-- (\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM9\ & ((\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM13\) # (\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM11\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000111111000000000011111100000011111111110000001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM11\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM13\,
	datad => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM9\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-11]_OTERM59\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-11]~4_combout\);

-- Location: FF_X19_Y61_N10
\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-12]_NEW_REG62\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~25_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-12]_OTERM63\);

-- Location: MLABCELL_X15_Y61_N9
\TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-12]~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-12]~3_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-12]_OTERM63\ & ( ((\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM13\ & 
-- \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM11\)) # (\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM9\) ) ) # ( !\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-12]_OTERM63\ & ( 
-- (\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM9\ & ((\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM11\) # (\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM13\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000011100000111000001110000011100011111000111110001111100011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM13\,
	datab => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM11\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM9\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-12]_OTERM63\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-12]~3_combout\);

-- Location: FF_X19_Y61_N8
\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-13]_NEW_REG90\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~21_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-13]_OTERM91\);

-- Location: MLABCELL_X15_Y61_N6
\TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-13]~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-13]~2_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-13]_OTERM91\ & ( ((\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM11\ & 
-- \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM13\)) # (\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM9\) ) ) # ( !\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-13]_OTERM91\ & ( 
-- (\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM9\ & ((\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM13\) # (\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM11\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000111111000000000011111100000011111111110000001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM11\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM13\,
	datad => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM9\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-13]_OTERM91\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-13]~2_combout\);

-- Location: FF_X19_Y61_N5
\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-14]_NEW_REG94\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~17_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-14]_OTERM95\);

-- Location: MLABCELL_X15_Y61_N33
\TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-14]~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-14]~1_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-14]_OTERM95\ & ( ((\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM13\ & 
-- \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM11\)) # (\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM9\) ) ) # ( !\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-14]_OTERM95\ & ( 
-- (\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM9\ & ((\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM11\) # (\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM13\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100001111000001010000111100001111010111110000111101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM13\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM9\,
	datad => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM11\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-14]_OTERM95\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-14]~1_combout\);

-- Location: FF_X19_Y61_N1
\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_NEW_REG14\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass1|Add3~13_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM15\);

-- Location: MLABCELL_X15_Y61_N15
\TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-15]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-15]~0_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM11\ & ( ((\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM15\ & 
-- \TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM13\)) # (\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM9\) ) ) # ( !\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM11\ & ( 
-- (\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM9\ & ((\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM13\) # (\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed[-15]_OTERM15\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000100110011001100110111011100010001001100110011001101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM15\,
	datab => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM9\,
	datad => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM13\,
	datae => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed[-15]_OTERM11\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-15]~0_combout\);

-- Location: MLABCELL_X15_Y62_N18
\TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-15]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-15]~0_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass1|Add4~5_sumout\ & ( (!\TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-15]~0_combout\ $ (!\TheRxFsk|Bandpasses:7:Bandpass1|Sum[-15]~q\)) # 
-- (\TheRxFsk|Bandpasses:7:Bandpass1|Add4~1_sumout\) ) ) # ( !\TheRxFsk|Bandpasses:7:Bandpass1|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:7:Bandpass1|Add4~1_sumout\ & (!\TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-15]~0_combout\ $ 
-- (!\TheRxFsk|Bandpasses:7:Bandpass1|Sum[-15]~q\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010101010000000001010101000001011111111101010101111111110101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~1_sumout\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResult[-15]~0_combout\,
	datad => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-15]~q\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~5_sumout\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-15]~0_combout\);

-- Location: FF_X15_Y62_N58
\TheRxFsk|Bandpasses:7:Bandpass1|R.SumState.SumEnable~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass1|Selector1~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass1|R.SumState.SumEnable~DUPLICATE_q\);

-- Location: LABCELL_X18_Y62_N54
\TheRxFsk|Bandpasses:7:Bandpass1|Selector2~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Selector2~0_combout\ = ((\TheRxFsk|Bandpasses:7:Bandpass1|R.SumState.SumSelect~q\ & ((!\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~0_combout\) # (!\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~1_combout\)))) # 
-- (\TheRxFsk|Bandpasses:7:Bandpass1|R.SumState.SumEnable~DUPLICATE_q\)

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111111101111000011111110111100001111111011110000111111101111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:11:Bandpass1|ALT_INV_Equal1~0_combout\,
	datab => \TheRxFsk|Bandpasses:11:Bandpass1|ALT_INV_Equal1~1_combout\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_R.SumState.SumEnable~DUPLICATE_q\,
	datad => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_R.SumState.SumSelect~q\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|Selector2~0_combout\);

-- Location: FF_X18_Y62_N55
\TheRxFsk|Bandpasses:7:Bandpass1|R.SumState.SumSelect\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass1|Selector2~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass1|R.SumState.SumSelect~q\);

-- Location: LABCELL_X18_Y62_N57
\TheRxFsk|Bandpasses:7:Bandpass1|Selector3~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Selector3~0_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass1|R.SumState.SumSelect~q\ & ( (\TheRxFsk|Bandpasses:11:Bandpass1|Equal1~0_combout\ & \TheRxFsk|Bandpasses:11:Bandpass1|Equal1~1_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000010001000100010001000100010001",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:11:Bandpass1|ALT_INV_Equal1~0_combout\,
	datab => \TheRxFsk|Bandpasses:11:Bandpass1|ALT_INV_Equal1~1_combout\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_R.SumState.SumSelect~q\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|Selector3~0_combout\);

-- Location: FF_X18_Y62_N59
\TheRxFsk|Bandpasses:7:Bandpass1|R.SumState.SumWait1\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass1|Selector3~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass1|R.SumState.SumWait1~q\);

-- Location: FF_X18_Y62_N4
\TheRxFsk|Bandpasses:7:Bandpass1|R.SumState.SumWait2\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	asdata => \TheRxFsk|Bandpasses:7:Bandpass1|R.SumState.SumWait1~q\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass1|R.SumState.SumWait2~q\);

-- Location: FF_X19_Y62_N40
\TheRxFsk|Bandpasses:7:Bandpass1|R.SumState.SumValid\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	asdata => \TheRxFsk|Bandpasses:7:Bandpass1|R.SumState.SumWait2~q\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass1|R.SumState.SumValid~q\);

-- Location: MLABCELL_X15_Y62_N15
\TheRxFsk|Bandpasses:7:Bandpass1|Selector0~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Selector0~0_combout\ = ( \TheI2sToPar|ValL~q\ & ( !\TheRxFsk|Bandpasses:7:Bandpass1|R.SumState.SumValid~q\ ) ) # ( !\TheI2sToPar|ValL~q\ & ( (!\TheRxFsk|Bandpasses:7:Bandpass1|R.SumState.SumValid~q\ & 
-- \TheRxFsk|Bandpasses:7:Bandpass1|R.SumState.Idle~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011110000000000001111000011110000111100001111000011110000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_R.SumState.SumValid~q\,
	datad => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_R.SumState.Idle~q\,
	dataf => \TheI2sToPar|ALT_INV_ValL~q\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|Selector0~0_combout\);

-- Location: FF_X15_Y62_N17
\TheRxFsk|Bandpasses:7:Bandpass1|R.SumState.Idle\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass1|Selector0~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass1|R.SumState.Idle~q\);

-- Location: MLABCELL_X15_Y62_N57
\TheRxFsk|Bandpasses:7:Bandpass1|Selector1~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Selector1~0_combout\ = ( \TheI2sToPar|ValL~q\ & ( !\TheRxFsk|Bandpasses:7:Bandpass1|R.SumState.Idle~q\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011110000111100001111000011110000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_R.SumState.Idle~q\,
	dataf => \TheI2sToPar|ALT_INV_ValL~q\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|Selector1~0_combout\);

-- Location: FF_X15_Y62_N59
\TheRxFsk|Bandpasses:7:Bandpass1|R.SumState.SumEnable\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass1|Selector1~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass1|R.SumState.SumEnable~q\);

-- Location: MLABCELL_X15_Y62_N12
\TheRxFsk|Bandpasses:7:Bandpass1|Selector6~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Selector6~0_combout\ = ((!\TheRxFsk|Bandpasses:7:Bandpass1|R.SumState.SumWait2~q\ & \TheRxFsk|Bandpasses:7:Bandpass1|R.SelSumUp~q\)) # (\TheRxFsk|Bandpasses:7:Bandpass1|R.SumState.SumEnable~q\)

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001111110011001100111111001100110011111100110011001111110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_R.SumState.SumEnable~q\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_R.SumState.SumWait2~q\,
	datad => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_R.SelSumUp~q\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|Selector6~0_combout\);

-- Location: FF_X15_Y62_N14
\TheRxFsk|Bandpasses:7:Bandpass1|R.SelSumUp\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass1|Selector6~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass1|R.SelSumUp~q\);

-- Location: MLABCELL_X15_Y62_N54
\TheRxFsk|Bandpasses:7:Bandpass1|Selector7~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Selector7~0_combout\ = ( \TheI2sToPar|ValL~q\ & ( (!\TheRxFsk|Bandpasses:7:Bandpass1|R.SumState.Idle~q\) # ((!\TheRxFsk|Bandpasses:7:Bandpass1|R.SumState.SumWait2~q\ & \TheRxFsk|Bandpasses:7:Bandpass1|R.EnableSumUp~q\)) ) 
-- ) # ( !\TheI2sToPar|ValL~q\ & ( (\TheRxFsk|Bandpasses:7:Bandpass1|R.EnableSumUp~q\ & ((!\TheRxFsk|Bandpasses:7:Bandpass1|R.SumState.SumWait2~q\) # (!\TheRxFsk|Bandpasses:7:Bandpass1|R.SumState.Idle~q\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011101110000000001110111011001100111011101100110011101110",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_R.SumState.SumWait2~q\,
	datab => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_R.SumState.Idle~q\,
	datad => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_R.EnableSumUp~q\,
	dataf => \TheI2sToPar|ALT_INV_ValL~q\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|Selector7~0_combout\);

-- Location: FF_X15_Y62_N56
\TheRxFsk|Bandpasses:7:Bandpass1|R.EnableSumUp\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass1|Selector7~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass1|R.EnableSumUp~q\);

-- Location: FF_X15_Y62_N19
\TheRxFsk|Bandpasses:7:Bandpass1|Sum[-15]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-15]~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:7:Bandpass1|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-15]~q\);

-- Location: LABCELL_X17_Y62_N0
\TheRxFsk|Bandpasses:7:Bandpass1|Add4~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add4~10\ = CARRY(( \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-15]~0_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-15]~q\ ) + ( !VCC ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000110011001100110000000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-15]~q\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResult[-15]~0_combout\,
	cin => GND,
	cout => \TheRxFsk|Bandpasses:7:Bandpass1|Add4~10\);

-- Location: LABCELL_X17_Y62_N3
\TheRxFsk|Bandpasses:7:Bandpass1|Add4~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add4~13_sumout\ = SUM(( \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-14]~1_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-14]~q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add4~10\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add4~14\ = CARRY(( \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-14]~1_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-14]~q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add4~10\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-14]~q\,
	datad => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResult[-14]~1_combout\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass1|Add4~10\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass1|Add4~13_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass1|Add4~14\);

-- Location: MLABCELL_X15_Y62_N3
\TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-14]~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-14]~1_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass1|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:7:Bandpass1|Add4~13_sumout\) # (\TheRxFsk|Bandpasses:7:Bandpass1|Add4~1_sumout\) ) ) # ( 
-- !\TheRxFsk|Bandpasses:7:Bandpass1|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:7:Bandpass1|Add4~1_sumout\ & \TheRxFsk|Bandpasses:7:Bandpass1|Add4~13_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100000101000001010000010101011111010111110101111101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~1_sumout\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~13_sumout\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~5_sumout\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-14]~1_combout\);

-- Location: FF_X15_Y62_N4
\TheRxFsk|Bandpasses:7:Bandpass1|Sum[-14]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-14]~1_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:7:Bandpass1|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-14]~q\);

-- Location: LABCELL_X17_Y62_N6
\TheRxFsk|Bandpasses:7:Bandpass1|Add4~17\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add4~17_sumout\ = SUM(( \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-13]~q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-13]~2_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add4~14\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add4~18\ = CARRY(( \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-13]~q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-13]~2_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add4~14\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111110000000000000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-13]~q\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResult[-13]~2_combout\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass1|Add4~14\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass1|Add4~17_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass1|Add4~18\);

-- Location: MLABCELL_X15_Y62_N24
\TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-13]~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-13]~2_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass1|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:7:Bandpass1|Add4~17_sumout\) # (\TheRxFsk|Bandpasses:7:Bandpass1|Add4~1_sumout\) ) ) # ( 
-- !\TheRxFsk|Bandpasses:7:Bandpass1|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:7:Bandpass1|Add4~1_sumout\ & \TheRxFsk|Bandpasses:7:Bandpass1|Add4~17_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100000101000001010000010101011111010111110101111101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~1_sumout\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~17_sumout\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~5_sumout\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-13]~2_combout\);

-- Location: FF_X15_Y62_N25
\TheRxFsk|Bandpasses:7:Bandpass1|Sum[-13]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-13]~2_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:7:Bandpass1|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-13]~q\);

-- Location: LABCELL_X17_Y62_N9
\TheRxFsk|Bandpasses:7:Bandpass1|Add4~21\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add4~21_sumout\ = SUM(( \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-12]~q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-12]~3_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add4~18\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add4~22\ = CARRY(( \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-12]~q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-12]~3_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add4~18\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000101010101010101000000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResult[-12]~3_combout\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-12]~q\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass1|Add4~18\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass1|Add4~21_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass1|Add4~22\);

-- Location: MLABCELL_X15_Y62_N27
\TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-12]~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-12]~3_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass1|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:7:Bandpass1|Add4~21_sumout\) # (\TheRxFsk|Bandpasses:7:Bandpass1|Add4~1_sumout\) ) ) # ( 
-- !\TheRxFsk|Bandpasses:7:Bandpass1|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:7:Bandpass1|Add4~1_sumout\ & \TheRxFsk|Bandpasses:7:Bandpass1|Add4~21_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100000101000001010000010101011111010111110101111101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~1_sumout\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~21_sumout\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~5_sumout\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-12]~3_combout\);

-- Location: FF_X15_Y62_N28
\TheRxFsk|Bandpasses:7:Bandpass1|Sum[-12]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-12]~3_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:7:Bandpass1|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-12]~q\);

-- Location: LABCELL_X17_Y62_N12
\TheRxFsk|Bandpasses:7:Bandpass1|Add4~25\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add4~25_sumout\ = SUM(( \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-11]~q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-11]~4_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add4~22\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add4~26\ = CARRY(( \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-11]~q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-11]~4_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add4~22\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-11]~q\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResult[-11]~4_combout\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass1|Add4~22\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass1|Add4~25_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass1|Add4~26\);

-- Location: MLABCELL_X15_Y62_N30
\TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-11]~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-11]~4_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass1|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:7:Bandpass1|Add4~25_sumout\) # (\TheRxFsk|Bandpasses:7:Bandpass1|Add4~1_sumout\) ) ) # ( 
-- !\TheRxFsk|Bandpasses:7:Bandpass1|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:7:Bandpass1|Add4~1_sumout\ & \TheRxFsk|Bandpasses:7:Bandpass1|Add4~25_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100000101000001010000010101011111010111110101111101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~1_sumout\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~25_sumout\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~5_sumout\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-11]~4_combout\);

-- Location: FF_X15_Y62_N31
\TheRxFsk|Bandpasses:7:Bandpass1|Sum[-11]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-11]~4_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:7:Bandpass1|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-11]~q\);

-- Location: LABCELL_X17_Y62_N15
\TheRxFsk|Bandpasses:7:Bandpass1|Add4~29\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add4~29_sumout\ = SUM(( \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-10]~q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-10]~5_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add4~26\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add4~30\ = CARRY(( \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-10]~q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-10]~5_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add4~26\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResult[-10]~5_combout\,
	datad => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-10]~q\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass1|Add4~26\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass1|Add4~29_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass1|Add4~30\);

-- Location: MLABCELL_X15_Y62_N33
\TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-10]~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-10]~5_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass1|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:7:Bandpass1|Add4~29_sumout\) # (\TheRxFsk|Bandpasses:7:Bandpass1|Add4~1_sumout\) ) ) # ( 
-- !\TheRxFsk|Bandpasses:7:Bandpass1|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:7:Bandpass1|Add4~1_sumout\ & \TheRxFsk|Bandpasses:7:Bandpass1|Add4~29_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100000101000001010000010101011111010111110101111101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~1_sumout\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~29_sumout\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~5_sumout\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-10]~5_combout\);

-- Location: FF_X15_Y62_N34
\TheRxFsk|Bandpasses:7:Bandpass1|Sum[-10]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-10]~5_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:7:Bandpass1|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-10]~q\);

-- Location: LABCELL_X17_Y62_N18
\TheRxFsk|Bandpasses:7:Bandpass1|Add4~33\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add4~33_sumout\ = SUM(( \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-9]~q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-9]~6_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add4~30\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add4~34\ = CARRY(( \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-9]~q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-9]~6_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add4~30\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000110011001100110000000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResult[-9]~6_combout\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-9]~q\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass1|Add4~30\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass1|Add4~33_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass1|Add4~34\);

-- Location: MLABCELL_X15_Y62_N36
\TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-9]~6\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-9]~6_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass1|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:7:Bandpass1|Add4~33_sumout\) # (\TheRxFsk|Bandpasses:7:Bandpass1|Add4~1_sumout\) ) ) # ( 
-- !\TheRxFsk|Bandpasses:7:Bandpass1|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:7:Bandpass1|Add4~1_sumout\ & \TheRxFsk|Bandpasses:7:Bandpass1|Add4~33_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100000101000001010000010101011111010111110101111101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~1_sumout\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~33_sumout\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~5_sumout\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-9]~6_combout\);

-- Location: FF_X15_Y62_N37
\TheRxFsk|Bandpasses:7:Bandpass1|Sum[-9]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-9]~6_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:7:Bandpass1|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-9]~q\);

-- Location: LABCELL_X17_Y62_N21
\TheRxFsk|Bandpasses:7:Bandpass1|Add4~37\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add4~37_sumout\ = SUM(( \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-8]~q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-8]~7_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add4~34\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add4~38\ = CARRY(( \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-8]~q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-8]~7_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add4~34\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-8]~q\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResult[-8]~7_combout\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass1|Add4~34\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass1|Add4~37_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass1|Add4~38\);

-- Location: MLABCELL_X15_Y62_N39
\TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-8]~7\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-8]~7_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass1|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:7:Bandpass1|Add4~37_sumout\) # (\TheRxFsk|Bandpasses:7:Bandpass1|Add4~1_sumout\) ) ) # ( 
-- !\TheRxFsk|Bandpasses:7:Bandpass1|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:7:Bandpass1|Add4~1_sumout\ & \TheRxFsk|Bandpasses:7:Bandpass1|Add4~37_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001010101000000000101010101010101111111110101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~1_sumout\,
	datad => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~37_sumout\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~5_sumout\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-8]~7_combout\);

-- Location: FF_X15_Y62_N40
\TheRxFsk|Bandpasses:7:Bandpass1|Sum[-8]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-8]~7_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:7:Bandpass1|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-8]~q\);

-- Location: LABCELL_X17_Y62_N24
\TheRxFsk|Bandpasses:7:Bandpass1|Add4~41\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add4~41_sumout\ = SUM(( \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-7]~q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-7]~8_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add4~38\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add4~42\ = CARRY(( \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-7]~q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-7]~8_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add4~38\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111110000000000000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-7]~q\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResult[-7]~8_combout\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass1|Add4~38\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass1|Add4~41_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass1|Add4~42\);

-- Location: MLABCELL_X15_Y62_N6
\TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-7]~8\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-7]~8_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass1|Add4~41_sumout\ & ( (\TheRxFsk|Bandpasses:7:Bandpass1|Add4~1_sumout\) # (\TheRxFsk|Bandpasses:7:Bandpass1|Add4~5_sumout\) ) ) # ( 
-- !\TheRxFsk|Bandpasses:7:Bandpass1|Add4~41_sumout\ & ( (\TheRxFsk|Bandpasses:7:Bandpass1|Add4~5_sumout\ & \TheRxFsk|Bandpasses:7:Bandpass1|Add4~1_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100000101000001010000010101011111010111110101111101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~5_sumout\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~1_sumout\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~41_sumout\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-7]~8_combout\);

-- Location: FF_X15_Y62_N7
\TheRxFsk|Bandpasses:7:Bandpass1|Sum[-7]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-7]~8_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:7:Bandpass1|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-7]~q\);

-- Location: LABCELL_X17_Y62_N27
\TheRxFsk|Bandpasses:7:Bandpass1|Add4~45\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add4~45_sumout\ = SUM(( \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-6]~q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-6]~9_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add4~42\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add4~46\ = CARRY(( \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-6]~q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-6]~9_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add4~42\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000110011001100110000000000000000000101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-6]~q\,
	datab => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResult[-6]~9_combout\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass1|Add4~42\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass1|Add4~45_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass1|Add4~46\);

-- Location: LABCELL_X16_Y62_N9
\TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-6]~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-6]~9_combout\ = (!\TheRxFsk|Bandpasses:7:Bandpass1|Add4~5_sumout\ & (\TheRxFsk|Bandpasses:7:Bandpass1|Add4~1_sumout\ & \TheRxFsk|Bandpasses:7:Bandpass1|Add4~45_sumout\)) # 
-- (\TheRxFsk|Bandpasses:7:Bandpass1|Add4~5_sumout\ & ((\TheRxFsk|Bandpasses:7:Bandpass1|Add4~45_sumout\) # (\TheRxFsk|Bandpasses:7:Bandpass1|Add4~1_sumout\)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010101011111000001010101111100000101010111110000010101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~5_sumout\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~1_sumout\,
	datad => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~45_sumout\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-6]~9_combout\);

-- Location: FF_X15_Y62_N11
\TheRxFsk|Bandpasses:7:Bandpass1|Sum[-6]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	asdata => \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-6]~9_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_R.SelSumUp~q\,
	sload => VCC,
	ena => \TheRxFsk|Bandpasses:7:Bandpass1|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-6]~q\);

-- Location: LABCELL_X17_Y62_N30
\TheRxFsk|Bandpasses:7:Bandpass1|Add4~49\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add4~49_sumout\ = SUM(( \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-5]~q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-5]~10_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add4~46\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add4~50\ = CARRY(( \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-5]~q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-5]~10_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add4~46\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-5]~q\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResult[-5]~10_combout\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass1|Add4~46\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass1|Add4~49_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass1|Add4~50\);

-- Location: MLABCELL_X15_Y62_N48
\TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-5]~10\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-5]~10_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass1|Add4~49_sumout\ & ( \TheRxFsk|Bandpasses:7:Bandpass1|Add4~5_sumout\ ) ) # ( !\TheRxFsk|Bandpasses:7:Bandpass1|Add4~49_sumout\ & ( 
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add4~5_sumout\ & ( \TheRxFsk|Bandpasses:7:Bandpass1|Add4~1_sumout\ ) ) ) # ( \TheRxFsk|Bandpasses:7:Bandpass1|Add4~49_sumout\ & ( !\TheRxFsk|Bandpasses:7:Bandpass1|Add4~5_sumout\ & ( 
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add4~1_sumout\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000011110000111100001111000011111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~1_sumout\,
	datae => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~49_sumout\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~5_sumout\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-5]~10_combout\);

-- Location: FF_X15_Y62_N49
\TheRxFsk|Bandpasses:7:Bandpass1|Sum[-5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-5]~10_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:7:Bandpass1|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-5]~q\);

-- Location: LABCELL_X17_Y62_N33
\TheRxFsk|Bandpasses:7:Bandpass1|Add4~53\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add4~53_sumout\ = SUM(( \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-4]~q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-4]~11_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add4~50\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add4~54\ = CARRY(( \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-4]~q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-4]~11_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add4~50\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111110000000000000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-4]~q\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResult[-4]~11_combout\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass1|Add4~50\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass1|Add4~53_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass1|Add4~54\);

-- Location: LABCELL_X16_Y62_N3
\TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-4]~11\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-4]~11_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass1|Add4~1_sumout\ & ( \TheRxFsk|Bandpasses:7:Bandpass1|Add4~5_sumout\ ) ) # ( !\TheRxFsk|Bandpasses:7:Bandpass1|Add4~1_sumout\ & ( 
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add4~5_sumout\ & ( \TheRxFsk|Bandpasses:7:Bandpass1|Add4~53_sumout\ ) ) ) # ( \TheRxFsk|Bandpasses:7:Bandpass1|Add4~1_sumout\ & ( !\TheRxFsk|Bandpasses:7:Bandpass1|Add4~5_sumout\ & ( 
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add4~53_sumout\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000010101010101010101010101010101011111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~53_sumout\,
	datae => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~1_sumout\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~5_sumout\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-4]~11_combout\);

-- Location: FF_X16_Y62_N4
\TheRxFsk|Bandpasses:7:Bandpass1|Sum[-4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-4]~11_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:7:Bandpass1|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-4]~q\);

-- Location: LABCELL_X17_Y62_N36
\TheRxFsk|Bandpasses:7:Bandpass1|Add4~57\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add4~57_sumout\ = SUM(( \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-3]~q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-3]~12_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add4~54\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add4~58\ = CARRY(( \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-3]~q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-3]~12_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add4~54\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000101010101010101000000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResult[-3]~12_combout\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-3]~q\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass1|Add4~54\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass1|Add4~57_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass1|Add4~58\);

-- Location: MLABCELL_X15_Y62_N42
\TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-3]~12\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-3]~12_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass1|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:7:Bandpass1|Add4~57_sumout\) # (\TheRxFsk|Bandpasses:7:Bandpass1|Add4~1_sumout\) ) ) # ( 
-- !\TheRxFsk|Bandpasses:7:Bandpass1|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:7:Bandpass1|Add4~1_sumout\ & \TheRxFsk|Bandpasses:7:Bandpass1|Add4~57_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000110011000000000011001100110011111111110011001111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~1_sumout\,
	datad => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~57_sumout\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~5_sumout\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-3]~12_combout\);

-- Location: FF_X15_Y62_N43
\TheRxFsk|Bandpasses:7:Bandpass1|Sum[-3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-3]~12_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:7:Bandpass1|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-3]~q\);

-- Location: LABCELL_X17_Y62_N39
\TheRxFsk|Bandpasses:7:Bandpass1|Add4~61\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add4~61_sumout\ = SUM(( \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-2]~q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-2]~13_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add4~58\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add4~62\ = CARRY(( \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-2]~q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-2]~13_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add4~58\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111110000000000000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-2]~q\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResult[-2]~13_combout\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass1|Add4~58\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass1|Add4~61_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass1|Add4~62\);

-- Location: MLABCELL_X15_Y62_N45
\TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-2]~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-2]~13_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass1|Add4~61_sumout\ & ( (\TheRxFsk|Bandpasses:7:Bandpass1|Add4~1_sumout\) # (\TheRxFsk|Bandpasses:7:Bandpass1|Add4~5_sumout\) ) ) # ( 
-- !\TheRxFsk|Bandpasses:7:Bandpass1|Add4~61_sumout\ & ( (\TheRxFsk|Bandpasses:7:Bandpass1|Add4~5_sumout\ & \TheRxFsk|Bandpasses:7:Bandpass1|Add4~1_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000100010001000100010001000101110111011101110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~5_sumout\,
	datab => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~1_sumout\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~61_sumout\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-2]~13_combout\);

-- Location: FF_X15_Y62_N46
\TheRxFsk|Bandpasses:7:Bandpass1|Sum[-2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-2]~13_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:7:Bandpass1|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-2]~q\);

-- Location: LABCELL_X17_Y62_N42
\TheRxFsk|Bandpasses:7:Bandpass1|Add4~65\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add4~65_sumout\ = SUM(( \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-1]~q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-1]~14_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add4~62\ ))
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add4~66\ = CARRY(( \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-1]~q\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|MultResult[-1]~14_combout\ ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add4~62\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000110011001100110000000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResult[-1]~14_combout\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-1]~q\,
	cin => \TheRxFsk|Bandpasses:7:Bandpass1|Add4~62\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass1|Add4~65_sumout\,
	cout => \TheRxFsk|Bandpasses:7:Bandpass1|Add4~66\);

-- Location: MLABCELL_X15_Y62_N21
\TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-1]~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-1]~14_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass1|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:7:Bandpass1|Add4~65_sumout\) # (\TheRxFsk|Bandpasses:7:Bandpass1|Add4~1_sumout\) ) ) # ( 
-- !\TheRxFsk|Bandpasses:7:Bandpass1|Add4~5_sumout\ & ( (\TheRxFsk|Bandpasses:7:Bandpass1|Add4~1_sumout\ & \TheRxFsk|Bandpasses:7:Bandpass1|Add4~65_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100000101000001010000010101011111010111110101111101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~1_sumout\,
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~65_sumout\,
	dataf => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~5_sumout\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-1]~14_combout\);

-- Location: FF_X15_Y62_N22
\TheRxFsk|Bandpasses:7:Bandpass1|Sum[-1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-1]~14_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:7:Bandpass1|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-1]~q\);

-- Location: LABCELL_X17_Y62_N48
\TheRxFsk|Bandpasses:7:Bandpass1|Add4~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add4~1_sumout\ = SUM(( \TheRxFsk|Bandpasses:7:Bandpass1|Sum\(0) ) + ( !\TheRxFsk|Bandpasses:7:Bandpass1|MultResultDelayed\(0) ) + ( \TheRxFsk|Bandpasses:7:Bandpass1|Add4~6\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000010101010101010100000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_MultResultDelayed\(0),
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum\(0),
	cin => \TheRxFsk|Bandpasses:7:Bandpass1|Add4~6\,
	sumout => \TheRxFsk|Bandpasses:7:Bandpass1|Add4~1_sumout\);

-- Location: MLABCELL_X15_Y62_N0
\TheRxFsk|Bandpasses:7:Bandpass1|Add4~1_wirecell\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Bandpasses:7:Bandpass1|Add4~1_wirecell_combout\ = !\TheRxFsk|Bandpasses:7:Bandpass1|Add4~1_sumout\

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1010101010101010101010101010101010101010101010101010101010101010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Add4~1_sumout\,
	combout => \TheRxFsk|Bandpasses:7:Bandpass1|Add4~1_wirecell_combout\);

-- Location: FF_X15_Y62_N1
\TheRxFsk|Bandpasses:7:Bandpass1|Sum[0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass1|Add4~1_wirecell_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:7:Bandpass1|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass1|Sum\(0));

-- Location: LABCELL_X24_Y60_N51
\TheRxFsk|Mux17~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Mux17~0_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-1]~q\ & ( (\TheRxFsk|Bandpasses:7:Bandpass1|Sum[-1]~q\) # (\SyncSwitchInput|Metastable\(1)) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass1|Sum[-1]~q\ & ( (!\SyncSwitchInput|Metastable\(1) & 
-- \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-1]~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000110000001100000011000000110000111111001111110011111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \SyncSwitchInput|ALT_INV_Metastable\(1),
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-1]~q\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-1]~q\,
	combout => \TheRxFsk|Mux17~0_combout\);

-- Location: LABCELL_X23_Y60_N18
\TheRxFsk|Mux18~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Mux18~0_combout\ = ( \SyncSwitchInput|Metastable\(1) & ( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-2]~q\ ) ) # ( !\SyncSwitchInput|Metastable\(1) & ( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-2]~q\ & ( \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-2]~q\ ) ) ) # 
-- ( !\SyncSwitchInput|Metastable\(1) & ( !\TheRxFsk|Bandpasses:4:Bandpass1|Sum[-2]~q\ & ( \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-2]~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111000000000000000000001111000011111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-2]~q\,
	datae => \SyncSwitchInput|ALT_INV_Metastable\(1),
	dataf => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-2]~q\,
	combout => \TheRxFsk|Mux18~0_combout\);

-- Location: FF_X15_Y62_N44
\TheRxFsk|Bandpasses:7:Bandpass1|Sum[-3]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Bandpasses:7:Bandpass1|NextSum[-3]~12_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Bandpasses:7:Bandpass1|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-3]~DUPLICATE_q\);

-- Location: LABCELL_X23_Y60_N15
\TheRxFsk|Mux19~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Mux19~0_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-3]~q\ & ( (\SyncSwitchInput|Metastable\(1)) # (\TheRxFsk|Bandpasses:7:Bandpass1|Sum[-3]~DUPLICATE_q\) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass1|Sum[-3]~q\ & ( 
-- (\TheRxFsk|Bandpasses:7:Bandpass1|Sum[-3]~DUPLICATE_q\ & !\SyncSwitchInput|Metastable\(1)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011000000110000001111110011111100110000001100000011111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-3]~DUPLICATE_q\,
	datac => \SyncSwitchInput|ALT_INV_Metastable\(1),
	datae => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-3]~q\,
	combout => \TheRxFsk|Mux19~0_combout\);

-- Location: LABCELL_X23_Y60_N57
\TheRxFsk|Mux20~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Mux20~0_combout\ = ( \SyncSwitchInput|Metastable\(1) & ( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-4]~q\ ) ) # ( !\SyncSwitchInput|Metastable\(1) & ( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-4]~q\ & ( \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-4]~q\ ) ) ) # 
-- ( !\SyncSwitchInput|Metastable\(1) & ( !\TheRxFsk|Bandpasses:4:Bandpass1|Sum[-4]~q\ & ( \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-4]~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111000000000000000000001111000011111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-4]~q\,
	datae => \SyncSwitchInput|ALT_INV_Metastable\(1),
	dataf => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-4]~q\,
	combout => \TheRxFsk|Mux20~0_combout\);

-- Location: MLABCELL_X21_Y64_N27
\TheRxFsk|Mux21~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Mux21~0_combout\ = ( \SyncSwitchInput|Metastable\(1) & ( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-5]~q\ ) ) # ( !\SyncSwitchInput|Metastable\(1) & ( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-5]~q\ & ( \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-5]~q\ ) ) ) # 
-- ( !\SyncSwitchInput|Metastable\(1) & ( !\TheRxFsk|Bandpasses:4:Bandpass1|Sum[-5]~q\ & ( \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-5]~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111000000000000000000001111000011111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-5]~q\,
	datae => \SyncSwitchInput|ALT_INV_Metastable\(1),
	dataf => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-5]~q\,
	combout => \TheRxFsk|Mux21~0_combout\);

-- Location: LABCELL_X23_Y60_N3
\TheRxFsk|Mux22~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Mux22~0_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-6]~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-6]~q\ ) ) # ( !\TheRxFsk|Bandpasses:7:Bandpass1|Sum[-6]~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-6]~q\ & ( 
-- \SyncSwitchInput|Metastable\(1) ) ) ) # ( \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-6]~q\ & ( !\TheRxFsk|Bandpasses:4:Bandpass1|Sum[-6]~q\ & ( !\SyncSwitchInput|Metastable\(1) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000001111000011111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \SyncSwitchInput|ALT_INV_Metastable\(1),
	datae => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-6]~q\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-6]~q\,
	combout => \TheRxFsk|Mux22~0_combout\);

-- Location: LABCELL_X23_Y60_N30
\TheRxFsk|Mux23~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Mux23~0_combout\ = ( \SyncSwitchInput|Metastable\(1) & ( \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-7]~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-7]~q\ ) ) ) # ( !\SyncSwitchInput|Metastable\(1) & ( \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-7]~q\ ) ) # 
-- ( \SyncSwitchInput|Metastable\(1) & ( !\TheRxFsk|Bandpasses:7:Bandpass1|Sum[-7]~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-7]~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000011110000111111111111111111110000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-7]~q\,
	datae => \SyncSwitchInput|ALT_INV_Metastable\(1),
	dataf => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-7]~q\,
	combout => \TheRxFsk|Mux23~0_combout\);

-- Location: LABCELL_X23_Y60_N51
\TheRxFsk|Mux24~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Mux24~0_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-8]~q\ & ( (!\SyncSwitchInput|Metastable\(1)) # (\TheRxFsk|Bandpasses:4:Bandpass1|Sum[-8]~q\) ) ) # ( !\TheRxFsk|Bandpasses:7:Bandpass1|Sum[-8]~q\ & ( 
-- (\TheRxFsk|Bandpasses:4:Bandpass1|Sum[-8]~q\ & \SyncSwitchInput|Metastable\(1)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100000011111100111111001100000011000000111111001111110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-8]~q\,
	datac => \SyncSwitchInput|ALT_INV_Metastable\(1),
	datae => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-8]~q\,
	combout => \TheRxFsk|Mux24~0_combout\);

-- Location: LABCELL_X23_Y60_N42
\TheRxFsk|Mux25~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Mux25~0_combout\ = ( \SyncSwitchInput|Metastable\(1) & ( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-9]~q\ ) ) # ( !\SyncSwitchInput|Metastable\(1) & ( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-9]~q\ & ( \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-9]~q\ ) ) ) # 
-- ( !\SyncSwitchInput|Metastable\(1) & ( !\TheRxFsk|Bandpasses:4:Bandpass1|Sum[-9]~q\ & ( \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-9]~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111000000000000000000001111000011111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-9]~q\,
	datae => \SyncSwitchInput|ALT_INV_Metastable\(1),
	dataf => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-9]~q\,
	combout => \TheRxFsk|Mux25~0_combout\);

-- Location: LABCELL_X24_Y60_N57
\TheRxFsk|Mux26~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Mux26~0_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-10]~q\ & ( (\TheRxFsk|Bandpasses:7:Bandpass1|Sum[-10]~q\) # (\SyncSwitchInput|Metastable\(1)) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass1|Sum[-10]~q\ & ( (!\SyncSwitchInput|Metastable\(1) 
-- & \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-10]~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000110000001100000011000000110000111111001111110011111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \SyncSwitchInput|ALT_INV_Metastable\(1),
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-10]~q\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-10]~q\,
	combout => \TheRxFsk|Mux26~0_combout\);

-- Location: LABCELL_X23_Y60_N36
\TheRxFsk|Mux27~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Mux27~0_combout\ = ( \SyncSwitchInput|Metastable\(1) & ( \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-11]~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-11]~q\ ) ) ) # ( !\SyncSwitchInput|Metastable\(1) & ( \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-11]~q\ ) 
-- ) # ( \SyncSwitchInput|Metastable\(1) & ( !\TheRxFsk|Bandpasses:7:Bandpass1|Sum[-11]~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-11]~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000001100110011001111111111111111110011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-11]~q\,
	datae => \SyncSwitchInput|ALT_INV_Metastable\(1),
	dataf => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-11]~q\,
	combout => \TheRxFsk|Mux27~0_combout\);

-- Location: LABCELL_X23_Y60_N6
\TheRxFsk|Mux28~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Mux28~0_combout\ = ( \SyncSwitchInput|Metastable\(1) & ( \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-12]~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-12]~q\ ) ) ) # ( !\SyncSwitchInput|Metastable\(1) & ( \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-12]~q\ ) 
-- ) # ( \SyncSwitchInput|Metastable\(1) & ( !\TheRxFsk|Bandpasses:7:Bandpass1|Sum[-12]~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-12]~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000011110000111111111111111111110000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-12]~q\,
	datae => \SyncSwitchInput|ALT_INV_Metastable\(1),
	dataf => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-12]~q\,
	combout => \TheRxFsk|Mux28~0_combout\);

-- Location: LABCELL_X23_Y60_N27
\TheRxFsk|Mux29~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Mux29~0_combout\ = ( \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-13]~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-13]~q\ ) ) # ( !\TheRxFsk|Bandpasses:7:Bandpass1|Sum[-13]~q\ & ( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-13]~q\ & ( 
-- \SyncSwitchInput|Metastable\(1) ) ) ) # ( \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-13]~q\ & ( !\TheRxFsk|Bandpasses:4:Bandpass1|Sum[-13]~q\ & ( !\SyncSwitchInput|Metastable\(1) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000001111000011111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \SyncSwitchInput|ALT_INV_Metastable\(1),
	datae => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-13]~q\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-13]~q\,
	combout => \TheRxFsk|Mux29~0_combout\);

-- Location: LABCELL_X24_Y60_N54
\TheRxFsk|Mux30~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Mux30~0_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-14]~q\ & ( (\TheRxFsk|Bandpasses:7:Bandpass1|Sum[-14]~q\) # (\SyncSwitchInput|Metastable\(1)) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass1|Sum[-14]~q\ & ( (!\SyncSwitchInput|Metastable\(1) 
-- & \TheRxFsk|Bandpasses:7:Bandpass1|Sum[-14]~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000110000001100000011000000110000111111001111110011111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \SyncSwitchInput|ALT_INV_Metastable\(1),
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-14]~q\,
	dataf => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-14]~q\,
	combout => \TheRxFsk|Mux30~0_combout\);

-- Location: LABCELL_X24_Y60_N48
\TheRxFsk|Mux31~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Mux31~0_combout\ = ( \TheRxFsk|Bandpasses:4:Bandpass1|Sum[-15]~q\ & ( (\SyncSwitchInput|Metastable\(1)) # (\TheRxFsk|Bandpasses:7:Bandpass1|Sum[-15]~q\) ) ) # ( !\TheRxFsk|Bandpasses:4:Bandpass1|Sum[-15]~q\ & ( 
-- (\TheRxFsk|Bandpasses:7:Bandpass1|Sum[-15]~q\ & !\SyncSwitchInput|Metastable\(1)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100000000000011110000000000001111111111110000111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum[-15]~q\,
	datad => \SyncSwitchInput|ALT_INV_Metastable\(1),
	dataf => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum[-15]~q\,
	combout => \TheRxFsk|Mux31~0_combout\);

-- Location: LABCELL_X24_Y60_N0
\TheRxFsk|Add1~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Add1~5_sumout\ = SUM(( (!\SyncSwitchInput|Metastable\(1) & (\TheRxFsk|Bandpasses:7:Bandpass1|Sum\(0))) # (\SyncSwitchInput|Metastable\(1) & ((\TheRxFsk|Bandpasses:4:Bandpass1|Sum\(0)))) ) + ( !\TheRxFsk|Mux31~0_combout\ $ 
-- (((!\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:7:Bandpass1|Sum\(0))) # (\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:4:Bandpass1|Sum\(0)))))) ) + ( !VCC ))
-- \TheRxFsk|Add1~6\ = CARRY(( (!\SyncSwitchInput|Metastable\(1) & (\TheRxFsk|Bandpasses:7:Bandpass1|Sum\(0))) # (\SyncSwitchInput|Metastable\(1) & ((\TheRxFsk|Bandpasses:4:Bandpass1|Sum\(0)))) ) + ( !\TheRxFsk|Mux31~0_combout\ $ 
-- (((!\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:7:Bandpass1|Sum\(0))) # (\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:4:Bandpass1|Sum\(0)))))) ) + ( !VCC ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000101110000100011100000000000000000100011101000111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum\(0),
	datab => \SyncSwitchInput|ALT_INV_Metastable\(1),
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum\(0),
	dataf => \TheRxFsk|ALT_INV_Mux31~0_combout\,
	cin => GND,
	sumout => \TheRxFsk|Add1~5_sumout\,
	cout => \TheRxFsk|Add1~6\);

-- Location: LABCELL_X24_Y60_N3
\TheRxFsk|Add1~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Add1~9_sumout\ = SUM(( !\TheRxFsk|Mux30~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:7:Bandpass1|Sum\(0))) # (\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:4:Bandpass1|Sum\(0)))))) ) + ( GND ) + ( 
-- \TheRxFsk|Add1~6\ ))
-- \TheRxFsk|Add1~10\ = CARRY(( !\TheRxFsk|Mux30~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:7:Bandpass1|Sum\(0))) # (\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:4:Bandpass1|Sum\(0)))))) ) + ( GND ) + ( 
-- \TheRxFsk|Add1~6\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000100011110111000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum\(0),
	datab => \SyncSwitchInput|ALT_INV_Metastable\(1),
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum\(0),
	datad => \TheRxFsk|ALT_INV_Mux30~0_combout\,
	cin => \TheRxFsk|Add1~6\,
	sumout => \TheRxFsk|Add1~9_sumout\,
	cout => \TheRxFsk|Add1~10\);

-- Location: LABCELL_X24_Y60_N6
\TheRxFsk|Add1~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Add1~13_sumout\ = SUM(( !\TheRxFsk|Mux29~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:7:Bandpass1|Sum\(0))) # (\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:4:Bandpass1|Sum\(0)))))) ) + ( GND ) + ( 
-- \TheRxFsk|Add1~10\ ))
-- \TheRxFsk|Add1~14\ = CARRY(( !\TheRxFsk|Mux29~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:7:Bandpass1|Sum\(0))) # (\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:4:Bandpass1|Sum\(0)))))) ) + ( GND ) + ( 
-- \TheRxFsk|Add1~10\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000100011110111000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum\(0),
	datab => \SyncSwitchInput|ALT_INV_Metastable\(1),
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum\(0),
	datad => \TheRxFsk|ALT_INV_Mux29~0_combout\,
	cin => \TheRxFsk|Add1~10\,
	sumout => \TheRxFsk|Add1~13_sumout\,
	cout => \TheRxFsk|Add1~14\);

-- Location: LABCELL_X24_Y60_N9
\TheRxFsk|Add1~17\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Add1~17_sumout\ = SUM(( !\TheRxFsk|Mux28~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:7:Bandpass1|Sum\(0))) # (\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:4:Bandpass1|Sum\(0)))))) ) + ( GND ) + ( 
-- \TheRxFsk|Add1~14\ ))
-- \TheRxFsk|Add1~18\ = CARRY(( !\TheRxFsk|Mux28~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:7:Bandpass1|Sum\(0))) # (\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:4:Bandpass1|Sum\(0)))))) ) + ( GND ) + ( 
-- \TheRxFsk|Add1~14\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000100011110111000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum\(0),
	datab => \SyncSwitchInput|ALT_INV_Metastable\(1),
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum\(0),
	datad => \TheRxFsk|ALT_INV_Mux28~0_combout\,
	cin => \TheRxFsk|Add1~14\,
	sumout => \TheRxFsk|Add1~17_sumout\,
	cout => \TheRxFsk|Add1~18\);

-- Location: LABCELL_X24_Y60_N12
\TheRxFsk|Add1~21\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Add1~21_sumout\ = SUM(( GND ) + ( !\TheRxFsk|Mux27~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:7:Bandpass1|Sum\(0))) # (\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:4:Bandpass1|Sum\(0)))))) ) + ( 
-- \TheRxFsk|Add1~18\ ))
-- \TheRxFsk|Add1~22\ = CARRY(( GND ) + ( !\TheRxFsk|Mux27~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:7:Bandpass1|Sum\(0))) # (\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:4:Bandpass1|Sum\(0)))))) ) + ( 
-- \TheRxFsk|Add1~18\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000101110000100011100000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum\(0),
	datab => \SyncSwitchInput|ALT_INV_Metastable\(1),
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum\(0),
	dataf => \TheRxFsk|ALT_INV_Mux27~0_combout\,
	cin => \TheRxFsk|Add1~18\,
	sumout => \TheRxFsk|Add1~21_sumout\,
	cout => \TheRxFsk|Add1~22\);

-- Location: LABCELL_X24_Y60_N15
\TheRxFsk|Add1~25\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Add1~25_sumout\ = SUM(( !\TheRxFsk|Mux26~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:7:Bandpass1|Sum\(0))) # (\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:4:Bandpass1|Sum\(0)))))) ) + ( GND ) + ( 
-- \TheRxFsk|Add1~22\ ))
-- \TheRxFsk|Add1~26\ = CARRY(( !\TheRxFsk|Mux26~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:7:Bandpass1|Sum\(0))) # (\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:4:Bandpass1|Sum\(0)))))) ) + ( GND ) + ( 
-- \TheRxFsk|Add1~22\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000100011110111000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum\(0),
	datab => \SyncSwitchInput|ALT_INV_Metastable\(1),
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum\(0),
	datad => \TheRxFsk|ALT_INV_Mux26~0_combout\,
	cin => \TheRxFsk|Add1~22\,
	sumout => \TheRxFsk|Add1~25_sumout\,
	cout => \TheRxFsk|Add1~26\);

-- Location: LABCELL_X24_Y60_N18
\TheRxFsk|Add1~29\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Add1~29_sumout\ = SUM(( !\TheRxFsk|Mux25~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:7:Bandpass1|Sum\(0))) # (\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:4:Bandpass1|Sum\(0)))))) ) + ( GND ) + ( 
-- \TheRxFsk|Add1~26\ ))
-- \TheRxFsk|Add1~30\ = CARRY(( !\TheRxFsk|Mux25~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:7:Bandpass1|Sum\(0))) # (\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:4:Bandpass1|Sum\(0)))))) ) + ( GND ) + ( 
-- \TheRxFsk|Add1~26\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000100011110111000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum\(0),
	datab => \SyncSwitchInput|ALT_INV_Metastable\(1),
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum\(0),
	datad => \TheRxFsk|ALT_INV_Mux25~0_combout\,
	cin => \TheRxFsk|Add1~26\,
	sumout => \TheRxFsk|Add1~29_sumout\,
	cout => \TheRxFsk|Add1~30\);

-- Location: LABCELL_X24_Y60_N21
\TheRxFsk|Add1~33\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Add1~33_sumout\ = SUM(( GND ) + ( !\TheRxFsk|Mux24~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:7:Bandpass1|Sum\(0))) # (\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:4:Bandpass1|Sum\(0)))))) ) + ( 
-- \TheRxFsk|Add1~30\ ))
-- \TheRxFsk|Add1~34\ = CARRY(( GND ) + ( !\TheRxFsk|Mux24~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:7:Bandpass1|Sum\(0))) # (\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:4:Bandpass1|Sum\(0)))))) ) + ( 
-- \TheRxFsk|Add1~30\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000101110000100011100000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum\(0),
	datab => \SyncSwitchInput|ALT_INV_Metastable\(1),
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum\(0),
	dataf => \TheRxFsk|ALT_INV_Mux24~0_combout\,
	cin => \TheRxFsk|Add1~30\,
	sumout => \TheRxFsk|Add1~33_sumout\,
	cout => \TheRxFsk|Add1~34\);

-- Location: LABCELL_X24_Y60_N24
\TheRxFsk|Add1~37\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Add1~37_sumout\ = SUM(( !\TheRxFsk|Mux23~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:7:Bandpass1|Sum\(0))) # (\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:4:Bandpass1|Sum\(0)))))) ) + ( GND ) + ( 
-- \TheRxFsk|Add1~34\ ))
-- \TheRxFsk|Add1~38\ = CARRY(( !\TheRxFsk|Mux23~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:7:Bandpass1|Sum\(0))) # (\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:4:Bandpass1|Sum\(0)))))) ) + ( GND ) + ( 
-- \TheRxFsk|Add1~34\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000100011110111000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum\(0),
	datab => \SyncSwitchInput|ALT_INV_Metastable\(1),
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum\(0),
	datad => \TheRxFsk|ALT_INV_Mux23~0_combout\,
	cin => \TheRxFsk|Add1~34\,
	sumout => \TheRxFsk|Add1~37_sumout\,
	cout => \TheRxFsk|Add1~38\);

-- Location: LABCELL_X24_Y60_N27
\TheRxFsk|Add1~41\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Add1~41_sumout\ = SUM(( GND ) + ( !\TheRxFsk|Mux22~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:7:Bandpass1|Sum\(0))) # (\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:4:Bandpass1|Sum\(0)))))) ) + ( 
-- \TheRxFsk|Add1~38\ ))
-- \TheRxFsk|Add1~42\ = CARRY(( GND ) + ( !\TheRxFsk|Mux22~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:7:Bandpass1|Sum\(0))) # (\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:4:Bandpass1|Sum\(0)))))) ) + ( 
-- \TheRxFsk|Add1~38\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000101110000100011100000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum\(0),
	datab => \SyncSwitchInput|ALT_INV_Metastable\(1),
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum\(0),
	dataf => \TheRxFsk|ALT_INV_Mux22~0_combout\,
	cin => \TheRxFsk|Add1~38\,
	sumout => \TheRxFsk|Add1~41_sumout\,
	cout => \TheRxFsk|Add1~42\);

-- Location: LABCELL_X24_Y60_N30
\TheRxFsk|Add1~45\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Add1~45_sumout\ = SUM(( !\TheRxFsk|Mux21~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:7:Bandpass1|Sum\(0))) # (\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:4:Bandpass1|Sum\(0)))))) ) + ( GND ) + ( 
-- \TheRxFsk|Add1~42\ ))
-- \TheRxFsk|Add1~46\ = CARRY(( !\TheRxFsk|Mux21~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:7:Bandpass1|Sum\(0))) # (\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:4:Bandpass1|Sum\(0)))))) ) + ( GND ) + ( 
-- \TheRxFsk|Add1~42\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000100011110111000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum\(0),
	datab => \SyncSwitchInput|ALT_INV_Metastable\(1),
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum\(0),
	datad => \TheRxFsk|ALT_INV_Mux21~0_combout\,
	cin => \TheRxFsk|Add1~42\,
	sumout => \TheRxFsk|Add1~45_sumout\,
	cout => \TheRxFsk|Add1~46\);

-- Location: LABCELL_X24_Y60_N33
\TheRxFsk|Add1~49\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Add1~49_sumout\ = SUM(( !\TheRxFsk|Mux20~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:7:Bandpass1|Sum\(0))) # (\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:4:Bandpass1|Sum\(0)))))) ) + ( GND ) + ( 
-- \TheRxFsk|Add1~46\ ))
-- \TheRxFsk|Add1~50\ = CARRY(( !\TheRxFsk|Mux20~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:7:Bandpass1|Sum\(0))) # (\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:4:Bandpass1|Sum\(0)))))) ) + ( GND ) + ( 
-- \TheRxFsk|Add1~46\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000100011110111000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum\(0),
	datab => \SyncSwitchInput|ALT_INV_Metastable\(1),
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum\(0),
	datad => \TheRxFsk|ALT_INV_Mux20~0_combout\,
	cin => \TheRxFsk|Add1~46\,
	sumout => \TheRxFsk|Add1~49_sumout\,
	cout => \TheRxFsk|Add1~50\);

-- Location: LABCELL_X24_Y60_N36
\TheRxFsk|Add1~53\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Add1~53_sumout\ = SUM(( GND ) + ( !\TheRxFsk|Mux19~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:7:Bandpass1|Sum\(0))) # (\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:4:Bandpass1|Sum\(0)))))) ) + ( 
-- \TheRxFsk|Add1~50\ ))
-- \TheRxFsk|Add1~54\ = CARRY(( GND ) + ( !\TheRxFsk|Mux19~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:7:Bandpass1|Sum\(0))) # (\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:4:Bandpass1|Sum\(0)))))) ) + ( 
-- \TheRxFsk|Add1~50\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000101110000100011100000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum\(0),
	datab => \SyncSwitchInput|ALT_INV_Metastable\(1),
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum\(0),
	dataf => \TheRxFsk|ALT_INV_Mux19~0_combout\,
	cin => \TheRxFsk|Add1~50\,
	sumout => \TheRxFsk|Add1~53_sumout\,
	cout => \TheRxFsk|Add1~54\);

-- Location: LABCELL_X24_Y60_N39
\TheRxFsk|Add1~57\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Add1~57_sumout\ = SUM(( GND ) + ( !\TheRxFsk|Mux18~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:7:Bandpass1|Sum\(0))) # (\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:4:Bandpass1|Sum\(0)))))) ) + ( 
-- \TheRxFsk|Add1~54\ ))
-- \TheRxFsk|Add1~58\ = CARRY(( GND ) + ( !\TheRxFsk|Mux18~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:7:Bandpass1|Sum\(0))) # (\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:4:Bandpass1|Sum\(0)))))) ) + ( 
-- \TheRxFsk|Add1~54\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000101110000100011100000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum\(0),
	datab => \SyncSwitchInput|ALT_INV_Metastable\(1),
	datac => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum\(0),
	dataf => \TheRxFsk|ALT_INV_Mux18~0_combout\,
	cin => \TheRxFsk|Add1~54\,
	sumout => \TheRxFsk|Add1~57_sumout\,
	cout => \TheRxFsk|Add1~58\);

-- Location: LABCELL_X24_Y60_N42
\TheRxFsk|Add1~61\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Add1~61_sumout\ = SUM(( GND ) + ( !\TheRxFsk|Mux17~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:7:Bandpass1|Sum\(0)))) # (\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:4:Bandpass1|Sum\(0))))) ) + ( 
-- \TheRxFsk|Add1~58\ ))
-- \TheRxFsk|Add1~62\ = CARRY(( GND ) + ( !\TheRxFsk|Mux17~0_combout\ $ (((!\SyncSwitchInput|Metastable\(1) & ((!\TheRxFsk|Bandpasses:7:Bandpass1|Sum\(0)))) # (\SyncSwitchInput|Metastable\(1) & (!\TheRxFsk|Bandpasses:4:Bandpass1|Sum\(0))))) ) + ( 
-- \TheRxFsk|Add1~58\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111000100001110100000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:4:Bandpass1|ALT_INV_Sum\(0),
	datab => \SyncSwitchInput|ALT_INV_Metastable\(1),
	datac => \TheRxFsk|Bandpasses:7:Bandpass1|ALT_INV_Sum\(0),
	dataf => \TheRxFsk|ALT_INV_Mux17~0_combout\,
	cin => \TheRxFsk|Add1~58\,
	sumout => \TheRxFsk|Add1~61_sumout\,
	cout => \TheRxFsk|Add1~62\);

-- Location: LABCELL_X24_Y60_N45
\TheRxFsk|Add1~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Add1~1_sumout\ = SUM(( GND ) + ( GND ) + ( \TheRxFsk|Add1~62\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	cin => \TheRxFsk|Add1~62\,
	sumout => \TheRxFsk|Add1~1_sumout\);

-- Location: LABCELL_X24_Y64_N0
\TheRxFsk|Add2~70\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Add2~70_cout\ = CARRY(( VCC ) + ( VCC ) + ( !VCC ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000000000001111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	cin => GND,
	cout => \TheRxFsk|Add2~70_cout\);

-- Location: LABCELL_X24_Y64_N3
\TheRxFsk|Add2~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Add2~9_sumout\ = SUM(( (\TheRxFsk|Add1~5_sumout\) # (\TheRxFsk|Add1~1_sumout\) ) + ( (!\TheRxFsk|Add0~1_sumout\ & !\TheRxFsk|Add0~5_sumout\) ) + ( \TheRxFsk|Add2~70_cout\ ))
-- \TheRxFsk|Add2~10\ = CARRY(( (\TheRxFsk|Add1~5_sumout\) # (\TheRxFsk|Add1~1_sumout\) ) + ( (!\TheRxFsk|Add0~1_sumout\ & !\TheRxFsk|Add0~5_sumout\) ) + ( \TheRxFsk|Add2~70_cout\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000010101011111111100000000000000000011111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|ALT_INV_Add0~1_sumout\,
	datab => \TheRxFsk|ALT_INV_Add1~1_sumout\,
	datac => \TheRxFsk|ALT_INV_Add1~5_sumout\,
	dataf => \TheRxFsk|ALT_INV_Add0~5_sumout\,
	cin => \TheRxFsk|Add2~70_cout\,
	sumout => \TheRxFsk|Add2~9_sumout\,
	cout => \TheRxFsk|Add2~10\);

-- Location: LABCELL_X24_Y64_N6
\TheRxFsk|Add2~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Add2~13_sumout\ = SUM(( (\TheRxFsk|Add1~9_sumout\) # (\TheRxFsk|Add1~1_sumout\) ) + ( (!\TheRxFsk|Add0~1_sumout\ & !\TheRxFsk|Add0~9_sumout\) ) + ( \TheRxFsk|Add2~10\ ))
-- \TheRxFsk|Add2~14\ = CARRY(( (\TheRxFsk|Add1~9_sumout\) # (\TheRxFsk|Add1~1_sumout\) ) + ( (!\TheRxFsk|Add0~1_sumout\ & !\TheRxFsk|Add0~9_sumout\) ) + ( \TheRxFsk|Add2~10\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000010101011111111100000000000000000011111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|ALT_INV_Add0~1_sumout\,
	datab => \TheRxFsk|ALT_INV_Add1~1_sumout\,
	datac => \TheRxFsk|ALT_INV_Add1~9_sumout\,
	dataf => \TheRxFsk|ALT_INV_Add0~9_sumout\,
	cin => \TheRxFsk|Add2~10\,
	sumout => \TheRxFsk|Add2~13_sumout\,
	cout => \TheRxFsk|Add2~14\);

-- Location: LABCELL_X24_Y64_N9
\TheRxFsk|Add2~17\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Add2~17_sumout\ = SUM(( (\TheRxFsk|Add1~13_sumout\) # (\TheRxFsk|Add1~1_sumout\) ) + ( (!\TheRxFsk|Add0~1_sumout\ & !\TheRxFsk|Add0~13_sumout\) ) + ( \TheRxFsk|Add2~14\ ))
-- \TheRxFsk|Add2~18\ = CARRY(( (\TheRxFsk|Add1~13_sumout\) # (\TheRxFsk|Add1~1_sumout\) ) + ( (!\TheRxFsk|Add0~1_sumout\ & !\TheRxFsk|Add0~13_sumout\) ) + ( \TheRxFsk|Add2~14\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000010101011111111100000000000000000011111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|ALT_INV_Add0~1_sumout\,
	datab => \TheRxFsk|ALT_INV_Add1~1_sumout\,
	datac => \TheRxFsk|ALT_INV_Add1~13_sumout\,
	dataf => \TheRxFsk|ALT_INV_Add0~13_sumout\,
	cin => \TheRxFsk|Add2~14\,
	sumout => \TheRxFsk|Add2~17_sumout\,
	cout => \TheRxFsk|Add2~18\);

-- Location: LABCELL_X24_Y64_N12
\TheRxFsk|Add2~21\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Add2~21_sumout\ = SUM(( (\TheRxFsk|Add1~17_sumout\) # (\TheRxFsk|Add1~1_sumout\) ) + ( (!\TheRxFsk|Add0~1_sumout\ & !\TheRxFsk|Add0~17_sumout\) ) + ( \TheRxFsk|Add2~18\ ))
-- \TheRxFsk|Add2~22\ = CARRY(( (\TheRxFsk|Add1~17_sumout\) # (\TheRxFsk|Add1~1_sumout\) ) + ( (!\TheRxFsk|Add0~1_sumout\ & !\TheRxFsk|Add0~17_sumout\) ) + ( \TheRxFsk|Add2~18\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000010101011111111100000000000000000011111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|ALT_INV_Add0~1_sumout\,
	datab => \TheRxFsk|ALT_INV_Add1~1_sumout\,
	datac => \TheRxFsk|ALT_INV_Add1~17_sumout\,
	dataf => \TheRxFsk|ALT_INV_Add0~17_sumout\,
	cin => \TheRxFsk|Add2~18\,
	sumout => \TheRxFsk|Add2~21_sumout\,
	cout => \TheRxFsk|Add2~22\);

-- Location: LABCELL_X24_Y64_N15
\TheRxFsk|Add2~25\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Add2~25_sumout\ = SUM(( (\TheRxFsk|Add1~21_sumout\) # (\TheRxFsk|Add1~1_sumout\) ) + ( (!\TheRxFsk|Add0~1_sumout\ & !\TheRxFsk|Add0~21_sumout\) ) + ( \TheRxFsk|Add2~22\ ))
-- \TheRxFsk|Add2~26\ = CARRY(( (\TheRxFsk|Add1~21_sumout\) # (\TheRxFsk|Add1~1_sumout\) ) + ( (!\TheRxFsk|Add0~1_sumout\ & !\TheRxFsk|Add0~21_sumout\) ) + ( \TheRxFsk|Add2~22\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000010101011111111100000000000000000011111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|ALT_INV_Add0~1_sumout\,
	datab => \TheRxFsk|ALT_INV_Add1~1_sumout\,
	datac => \TheRxFsk|ALT_INV_Add1~21_sumout\,
	dataf => \TheRxFsk|ALT_INV_Add0~21_sumout\,
	cin => \TheRxFsk|Add2~22\,
	sumout => \TheRxFsk|Add2~25_sumout\,
	cout => \TheRxFsk|Add2~26\);

-- Location: LABCELL_X24_Y64_N18
\TheRxFsk|Add2~29\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Add2~29_sumout\ = SUM(( (\TheRxFsk|Add1~25_sumout\) # (\TheRxFsk|Add1~1_sumout\) ) + ( (!\TheRxFsk|Add0~1_sumout\ & !\TheRxFsk|Add0~25_sumout\) ) + ( \TheRxFsk|Add2~26\ ))
-- \TheRxFsk|Add2~30\ = CARRY(( (\TheRxFsk|Add1~25_sumout\) # (\TheRxFsk|Add1~1_sumout\) ) + ( (!\TheRxFsk|Add0~1_sumout\ & !\TheRxFsk|Add0~25_sumout\) ) + ( \TheRxFsk|Add2~26\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000010101011111111100000000000000000011111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|ALT_INV_Add0~1_sumout\,
	datab => \TheRxFsk|ALT_INV_Add1~1_sumout\,
	datac => \TheRxFsk|ALT_INV_Add1~25_sumout\,
	dataf => \TheRxFsk|ALT_INV_Add0~25_sumout\,
	cin => \TheRxFsk|Add2~26\,
	sumout => \TheRxFsk|Add2~29_sumout\,
	cout => \TheRxFsk|Add2~30\);

-- Location: LABCELL_X24_Y64_N21
\TheRxFsk|Add2~33\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Add2~33_sumout\ = SUM(( (\TheRxFsk|Add1~29_sumout\) # (\TheRxFsk|Add1~1_sumout\) ) + ( (!\TheRxFsk|Add0~1_sumout\ & !\TheRxFsk|Add0~29_sumout\) ) + ( \TheRxFsk|Add2~30\ ))
-- \TheRxFsk|Add2~34\ = CARRY(( (\TheRxFsk|Add1~29_sumout\) # (\TheRxFsk|Add1~1_sumout\) ) + ( (!\TheRxFsk|Add0~1_sumout\ & !\TheRxFsk|Add0~29_sumout\) ) + ( \TheRxFsk|Add2~30\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000010101011111111100000000000000000011111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|ALT_INV_Add0~1_sumout\,
	datab => \TheRxFsk|ALT_INV_Add1~1_sumout\,
	datac => \TheRxFsk|ALT_INV_Add1~29_sumout\,
	dataf => \TheRxFsk|ALT_INV_Add0~29_sumout\,
	cin => \TheRxFsk|Add2~30\,
	sumout => \TheRxFsk|Add2~33_sumout\,
	cout => \TheRxFsk|Add2~34\);

-- Location: LABCELL_X24_Y64_N24
\TheRxFsk|Add2~37\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Add2~37_sumout\ = SUM(( (\TheRxFsk|Add1~33_sumout\) # (\TheRxFsk|Add1~1_sumout\) ) + ( (!\TheRxFsk|Add0~1_sumout\ & !\TheRxFsk|Add0~33_sumout\) ) + ( \TheRxFsk|Add2~34\ ))
-- \TheRxFsk|Add2~38\ = CARRY(( (\TheRxFsk|Add1~33_sumout\) # (\TheRxFsk|Add1~1_sumout\) ) + ( (!\TheRxFsk|Add0~1_sumout\ & !\TheRxFsk|Add0~33_sumout\) ) + ( \TheRxFsk|Add2~34\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000010101011111111100000000000000000011111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|ALT_INV_Add0~1_sumout\,
	datab => \TheRxFsk|ALT_INV_Add1~1_sumout\,
	datac => \TheRxFsk|ALT_INV_Add1~33_sumout\,
	dataf => \TheRxFsk|ALT_INV_Add0~33_sumout\,
	cin => \TheRxFsk|Add2~34\,
	sumout => \TheRxFsk|Add2~37_sumout\,
	cout => \TheRxFsk|Add2~38\);

-- Location: LABCELL_X24_Y64_N27
\TheRxFsk|Add2~41\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Add2~41_sumout\ = SUM(( (\TheRxFsk|Add1~37_sumout\) # (\TheRxFsk|Add1~1_sumout\) ) + ( (!\TheRxFsk|Add0~1_sumout\ & !\TheRxFsk|Add0~37_sumout\) ) + ( \TheRxFsk|Add2~38\ ))
-- \TheRxFsk|Add2~42\ = CARRY(( (\TheRxFsk|Add1~37_sumout\) # (\TheRxFsk|Add1~1_sumout\) ) + ( (!\TheRxFsk|Add0~1_sumout\ & !\TheRxFsk|Add0~37_sumout\) ) + ( \TheRxFsk|Add2~38\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000010101011111111100000000000000000011111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|ALT_INV_Add0~1_sumout\,
	datab => \TheRxFsk|ALT_INV_Add1~1_sumout\,
	datac => \TheRxFsk|ALT_INV_Add1~37_sumout\,
	dataf => \TheRxFsk|ALT_INV_Add0~37_sumout\,
	cin => \TheRxFsk|Add2~38\,
	sumout => \TheRxFsk|Add2~41_sumout\,
	cout => \TheRxFsk|Add2~42\);

-- Location: LABCELL_X24_Y64_N30
\TheRxFsk|Add2~45\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Add2~45_sumout\ = SUM(( (!\TheRxFsk|Add0~1_sumout\ & !\TheRxFsk|Add0~41_sumout\) ) + ( (\TheRxFsk|Add1~41_sumout\) # (\TheRxFsk|Add1~1_sumout\) ) + ( \TheRxFsk|Add2~42\ ))
-- \TheRxFsk|Add2~46\ = CARRY(( (!\TheRxFsk|Add0~1_sumout\ & !\TheRxFsk|Add0~41_sumout\) ) + ( (\TheRxFsk|Add1~41_sumout\) # (\TheRxFsk|Add1~1_sumout\) ) + ( \TheRxFsk|Add2~42\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000110011000000000000000000000000001010000010100000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|ALT_INV_Add0~1_sumout\,
	datab => \TheRxFsk|ALT_INV_Add1~1_sumout\,
	datac => \TheRxFsk|ALT_INV_Add0~41_sumout\,
	dataf => \TheRxFsk|ALT_INV_Add1~41_sumout\,
	cin => \TheRxFsk|Add2~42\,
	sumout => \TheRxFsk|Add2~45_sumout\,
	cout => \TheRxFsk|Add2~46\);

-- Location: LABCELL_X24_Y64_N33
\TheRxFsk|Add2~49\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Add2~49_sumout\ = SUM(( (\TheRxFsk|Add1~45_sumout\) # (\TheRxFsk|Add1~1_sumout\) ) + ( (!\TheRxFsk|Add0~1_sumout\ & !\TheRxFsk|Add0~45_sumout\) ) + ( \TheRxFsk|Add2~46\ ))
-- \TheRxFsk|Add2~50\ = CARRY(( (\TheRxFsk|Add1~45_sumout\) # (\TheRxFsk|Add1~1_sumout\) ) + ( (!\TheRxFsk|Add0~1_sumout\ & !\TheRxFsk|Add0~45_sumout\) ) + ( \TheRxFsk|Add2~46\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000010101011111111100000000000000000011111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|ALT_INV_Add0~1_sumout\,
	datab => \TheRxFsk|ALT_INV_Add1~1_sumout\,
	datac => \TheRxFsk|ALT_INV_Add1~45_sumout\,
	dataf => \TheRxFsk|ALT_INV_Add0~45_sumout\,
	cin => \TheRxFsk|Add2~46\,
	sumout => \TheRxFsk|Add2~49_sumout\,
	cout => \TheRxFsk|Add2~50\);

-- Location: LABCELL_X24_Y64_N36
\TheRxFsk|Add2~53\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Add2~53_sumout\ = SUM(( (\TheRxFsk|Add1~49_sumout\) # (\TheRxFsk|Add1~1_sumout\) ) + ( (!\TheRxFsk|Add0~1_sumout\ & !\TheRxFsk|Add0~49_sumout\) ) + ( \TheRxFsk|Add2~50\ ))
-- \TheRxFsk|Add2~54\ = CARRY(( (\TheRxFsk|Add1~49_sumout\) # (\TheRxFsk|Add1~1_sumout\) ) + ( (!\TheRxFsk|Add0~1_sumout\ & !\TheRxFsk|Add0~49_sumout\) ) + ( \TheRxFsk|Add2~50\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000010101011111111100000000000000000011111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|ALT_INV_Add0~1_sumout\,
	datab => \TheRxFsk|ALT_INV_Add1~1_sumout\,
	datac => \TheRxFsk|ALT_INV_Add1~49_sumout\,
	dataf => \TheRxFsk|ALT_INV_Add0~49_sumout\,
	cin => \TheRxFsk|Add2~50\,
	sumout => \TheRxFsk|Add2~53_sumout\,
	cout => \TheRxFsk|Add2~54\);

-- Location: LABCELL_X24_Y64_N39
\TheRxFsk|Add2~57\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Add2~57_sumout\ = SUM(( (!\TheRxFsk|Add0~1_sumout\ & !\TheRxFsk|Add0~53_sumout\) ) + ( (\TheRxFsk|Add1~53_sumout\) # (\TheRxFsk|Add1~1_sumout\) ) + ( \TheRxFsk|Add2~54\ ))
-- \TheRxFsk|Add2~58\ = CARRY(( (!\TheRxFsk|Add0~1_sumout\ & !\TheRxFsk|Add0~53_sumout\) ) + ( (\TheRxFsk|Add1~53_sumout\) # (\TheRxFsk|Add1~1_sumout\) ) + ( \TheRxFsk|Add2~54\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000110011000000000000000000000000001010000010100000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|ALT_INV_Add0~1_sumout\,
	datab => \TheRxFsk|ALT_INV_Add1~1_sumout\,
	datac => \TheRxFsk|ALT_INV_Add0~53_sumout\,
	dataf => \TheRxFsk|ALT_INV_Add1~53_sumout\,
	cin => \TheRxFsk|Add2~54\,
	sumout => \TheRxFsk|Add2~57_sumout\,
	cout => \TheRxFsk|Add2~58\);

-- Location: LABCELL_X24_Y64_N42
\TheRxFsk|Add2~61\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Add2~61_sumout\ = SUM(( (\TheRxFsk|Add1~57_sumout\) # (\TheRxFsk|Add1~1_sumout\) ) + ( (!\TheRxFsk|Add0~1_sumout\ & !\TheRxFsk|Add0~57_sumout\) ) + ( \TheRxFsk|Add2~58\ ))
-- \TheRxFsk|Add2~62\ = CARRY(( (\TheRxFsk|Add1~57_sumout\) # (\TheRxFsk|Add1~1_sumout\) ) + ( (!\TheRxFsk|Add0~1_sumout\ & !\TheRxFsk|Add0~57_sumout\) ) + ( \TheRxFsk|Add2~58\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000010101011111111100000000000000000011111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|ALT_INV_Add0~1_sumout\,
	datab => \TheRxFsk|ALT_INV_Add1~1_sumout\,
	datac => \TheRxFsk|ALT_INV_Add1~57_sumout\,
	dataf => \TheRxFsk|ALT_INV_Add0~57_sumout\,
	cin => \TheRxFsk|Add2~58\,
	sumout => \TheRxFsk|Add2~61_sumout\,
	cout => \TheRxFsk|Add2~62\);

-- Location: LABCELL_X24_Y64_N45
\TheRxFsk|Add2~65\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Add2~65_sumout\ = SUM(( (!\TheRxFsk|Add0~1_sumout\ & !\TheRxFsk|Add0~61_sumout\) ) + ( (\TheRxFsk|Add1~61_sumout\) # (\TheRxFsk|Add1~1_sumout\) ) + ( \TheRxFsk|Add2~62\ ))
-- \TheRxFsk|Add2~66\ = CARRY(( (!\TheRxFsk|Add0~1_sumout\ & !\TheRxFsk|Add0~61_sumout\) ) + ( (\TheRxFsk|Add1~61_sumout\) # (\TheRxFsk|Add1~1_sumout\) ) + ( \TheRxFsk|Add2~62\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000110011000000000000000000000000001010000010100000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|ALT_INV_Add0~1_sumout\,
	datab => \TheRxFsk|ALT_INV_Add1~1_sumout\,
	datac => \TheRxFsk|ALT_INV_Add0~61_sumout\,
	dataf => \TheRxFsk|ALT_INV_Add1~61_sumout\,
	cin => \TheRxFsk|Add2~62\,
	sumout => \TheRxFsk|Add2~65_sumout\,
	cout => \TheRxFsk|Add2~66\);

-- Location: LABCELL_X24_Y64_N48
\TheRxFsk|Add2~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Add2~1_sumout\ = SUM(( VCC ) + ( GND ) + ( \TheRxFsk|Add2~66\ ))
-- \TheRxFsk|Add2~2\ = CARRY(( VCC ) + ( GND ) + ( \TheRxFsk|Add2~66\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000001111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	cin => \TheRxFsk|Add2~66\,
	sumout => \TheRxFsk|Add2~1_sumout\,
	cout => \TheRxFsk|Add2~2\);

-- Location: LABCELL_X24_Y64_N51
\TheRxFsk|Add2~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Add2~5_sumout\ = SUM(( VCC ) + ( GND ) + ( \TheRxFsk|Add2~2\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000001111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	cin => \TheRxFsk|Add2~2\,
	sumout => \TheRxFsk|Add2~5_sumout\);

-- Location: MLABCELL_X25_Y64_N27
\TheRxFsk|Substracted[-15]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Substracted[-15]~0_combout\ = ( \TheRxFsk|Add2~9_sumout\ & ( (!\TheRxFsk|Add2~5_sumout\) # (\TheRxFsk|Add2~1_sumout\) ) ) # ( !\TheRxFsk|Add2~9_sumout\ & ( (!\TheRxFsk|Add2~5_sumout\ & \TheRxFsk|Add2~1_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000101000001010000010100000101010101111101011111010111110101111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|ALT_INV_Add2~5_sumout\,
	datac => \TheRxFsk|ALT_INV_Add2~1_sumout\,
	dataf => \TheRxFsk|ALT_INV_Add2~9_sumout\,
	combout => \TheRxFsk|Substracted[-15]~0_combout\);

-- Location: MLABCELL_X28_Y64_N27
\TheRxFsk|Lowpass|R.WriteAddress[0]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|R.WriteAddress[0]~0_combout\ = ( \TheRxFsk|Lowpass|CoefMemory~0_combout\ & ( (\TheRxFsk|Lowpass|Equal1~0_combout\ & \TheRxFsk|Lowpass|R.AddressState~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000000011110000000000001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Lowpass|ALT_INV_Equal1~0_combout\,
	datad => \TheRxFsk|Lowpass|ALT_INV_R.AddressState~q\,
	dataf => \TheRxFsk|Lowpass|ALT_INV_CoefMemory~0_combout\,
	combout => \TheRxFsk|Lowpass|R.WriteAddress[0]~0_combout\);

-- Location: FF_X27_Y64_N26
\TheRxFsk|Lowpass|R.WriteAddress[0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|vNextWriteAddress~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	ena => \TheRxFsk|Lowpass|R.WriteAddress[0]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|R.WriteAddress\(0));

-- Location: LABCELL_X27_Y64_N0
\TheRxFsk|Lowpass|Add1~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add1~2\ = CARRY(( \TheRxFsk|Lowpass|R.WriteAddress\(0) ) + ( VCC ) + ( !VCC ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Lowpass|ALT_INV_R.WriteAddress\(0),
	cin => GND,
	cout => \TheRxFsk|Lowpass|Add1~2\);

-- Location: LABCELL_X27_Y64_N3
\TheRxFsk|Lowpass|Add1~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add1~5_sumout\ = SUM(( !\TheRxFsk|Lowpass|R.WriteAddress\(1) ) + ( VCC ) + ( \TheRxFsk|Lowpass|Add1~2\ ))
-- \TheRxFsk|Lowpass|Add1~6\ = CARRY(( !\TheRxFsk|Lowpass|R.WriteAddress\(1) ) + ( VCC ) + ( \TheRxFsk|Lowpass|Add1~2\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000000000001111000011110000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Lowpass|ALT_INV_R.WriteAddress\(1),
	cin => \TheRxFsk|Lowpass|Add1~2\,
	sumout => \TheRxFsk|Lowpass|Add1~5_sumout\,
	cout => \TheRxFsk|Lowpass|Add1~6\);

-- Location: LABCELL_X27_Y64_N42
\TheRxFsk|Lowpass|R.WriteAddress[1]~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|R.WriteAddress[1]~1_combout\ = !\TheRxFsk|Lowpass|Add1~5_sumout\

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111000011110000111100001111000011110000111100001111000011110000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Lowpass|ALT_INV_Add1~5_sumout\,
	combout => \TheRxFsk|Lowpass|R.WriteAddress[1]~1_combout\);

-- Location: FF_X27_Y64_N44
\TheRxFsk|Lowpass|R.WriteAddress[1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|R.WriteAddress[1]~1_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	ena => \TheRxFsk|Lowpass|R.WriteAddress[0]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|R.WriteAddress\(1));

-- Location: LABCELL_X27_Y64_N6
\TheRxFsk|Lowpass|Add1~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add1~9_sumout\ = SUM(( \TheRxFsk|Lowpass|R.WriteAddress\(2) ) + ( VCC ) + ( \TheRxFsk|Lowpass|Add1~6\ ))
-- \TheRxFsk|Lowpass|Add1~10\ = CARRY(( \TheRxFsk|Lowpass|R.WriteAddress\(2) ) + ( VCC ) + ( \TheRxFsk|Lowpass|Add1~6\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Lowpass|ALT_INV_R.WriteAddress\(2),
	cin => \TheRxFsk|Lowpass|Add1~6\,
	sumout => \TheRxFsk|Lowpass|Add1~9_sumout\,
	cout => \TheRxFsk|Lowpass|Add1~10\);

-- Location: LABCELL_X27_Y64_N48
\TheRxFsk|Lowpass|vNextWriteAddress~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|vNextWriteAddress~1_combout\ = ( \TheRxFsk|Lowpass|Add1~9_sumout\ & ( ((!\TheRxFsk|Lowpass|R.WriteAddress\(1)) # ((!\TheRxFsk|Lowpass|Equal2~0_combout\) # (\TheRxFsk|Lowpass|R.WriteAddress\(2)))) # (\TheRxFsk|Lowpass|R.WriteAddress\(0)) 
-- ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111101111111111111110111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_R.WriteAddress\(0),
	datab => \TheRxFsk|Lowpass|ALT_INV_R.WriteAddress\(1),
	datac => \TheRxFsk|Lowpass|ALT_INV_Equal2~0_combout\,
	datad => \TheRxFsk|Lowpass|ALT_INV_R.WriteAddress\(2),
	dataf => \TheRxFsk|Lowpass|ALT_INV_Add1~9_sumout\,
	combout => \TheRxFsk|Lowpass|vNextWriteAddress~1_combout\);

-- Location: FF_X27_Y64_N50
\TheRxFsk|Lowpass|R.WriteAddress[2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|vNextWriteAddress~1_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	ena => \TheRxFsk|Lowpass|R.WriteAddress[0]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|R.WriteAddress\(2));

-- Location: LABCELL_X27_Y64_N9
\TheRxFsk|Lowpass|Add1~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add1~13_sumout\ = SUM(( !\TheRxFsk|Lowpass|R.WriteAddress\(3) ) + ( VCC ) + ( \TheRxFsk|Lowpass|Add1~10\ ))
-- \TheRxFsk|Lowpass|Add1~14\ = CARRY(( !\TheRxFsk|Lowpass|R.WriteAddress\(3) ) + ( VCC ) + ( \TheRxFsk|Lowpass|Add1~10\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000000000001111000011110000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Lowpass|ALT_INV_R.WriteAddress\(3),
	cin => \TheRxFsk|Lowpass|Add1~10\,
	sumout => \TheRxFsk|Lowpass|Add1~13_sumout\,
	cout => \TheRxFsk|Lowpass|Add1~14\);

-- Location: LABCELL_X27_Y64_N45
\TheRxFsk|Lowpass|R.WriteAddress[3]~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|R.WriteAddress[3]~2_combout\ = ( !\TheRxFsk|Lowpass|Add1~13_sumout\ )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111111111111111111111111111100000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \TheRxFsk|Lowpass|ALT_INV_Add1~13_sumout\,
	combout => \TheRxFsk|Lowpass|R.WriteAddress[3]~2_combout\);

-- Location: FF_X27_Y64_N47
\TheRxFsk|Lowpass|R.WriteAddress[3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|R.WriteAddress[3]~2_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	ena => \TheRxFsk|Lowpass|R.WriteAddress[0]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|R.WriteAddress\(3));

-- Location: LABCELL_X27_Y64_N12
\TheRxFsk|Lowpass|Add1~17\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add1~17_sumout\ = SUM(( \TheRxFsk|Lowpass|R.WriteAddress\(4) ) + ( VCC ) + ( \TheRxFsk|Lowpass|Add1~14\ ))
-- \TheRxFsk|Lowpass|Add1~18\ = CARRY(( \TheRxFsk|Lowpass|R.WriteAddress\(4) ) + ( VCC ) + ( \TheRxFsk|Lowpass|Add1~14\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000000000000011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Lowpass|ALT_INV_R.WriteAddress\(4),
	cin => \TheRxFsk|Lowpass|Add1~14\,
	sumout => \TheRxFsk|Lowpass|Add1~17_sumout\,
	cout => \TheRxFsk|Lowpass|Add1~18\);

-- Location: LABCELL_X27_Y64_N51
\TheRxFsk|Lowpass|vNextWriteAddress~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|vNextWriteAddress~2_combout\ = ( \TheRxFsk|Lowpass|R.WriteAddress\(2) & ( \TheRxFsk|Lowpass|Add1~17_sumout\ ) ) # ( !\TheRxFsk|Lowpass|R.WriteAddress\(2) & ( (\TheRxFsk|Lowpass|Add1~17_sumout\ & (((!\TheRxFsk|Lowpass|R.WriteAddress\(1)) 
-- # (!\TheRxFsk|Lowpass|Equal2~0_combout\)) # (\TheRxFsk|Lowpass|R.WriteAddress\(0)))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001101000011110000110100001111000011110000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_R.WriteAddress\(0),
	datab => \TheRxFsk|Lowpass|ALT_INV_R.WriteAddress\(1),
	datac => \TheRxFsk|Lowpass|ALT_INV_Add1~17_sumout\,
	datad => \TheRxFsk|Lowpass|ALT_INV_Equal2~0_combout\,
	dataf => \TheRxFsk|Lowpass|ALT_INV_R.WriteAddress\(2),
	combout => \TheRxFsk|Lowpass|vNextWriteAddress~2_combout\);

-- Location: FF_X27_Y64_N52
\TheRxFsk|Lowpass|R.WriteAddress[4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|vNextWriteAddress~2_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	ena => \TheRxFsk|Lowpass|R.WriteAddress[0]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|R.WriteAddress\(4));

-- Location: LABCELL_X27_Y64_N15
\TheRxFsk|Lowpass|Add1~21\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add1~21_sumout\ = SUM(( \TheRxFsk|Lowpass|R.WriteAddress\(5) ) + ( VCC ) + ( \TheRxFsk|Lowpass|Add1~18\ ))
-- \TheRxFsk|Lowpass|Add1~22\ = CARRY(( \TheRxFsk|Lowpass|R.WriteAddress\(5) ) + ( VCC ) + ( \TheRxFsk|Lowpass|Add1~18\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Lowpass|ALT_INV_R.WriteAddress\(5),
	cin => \TheRxFsk|Lowpass|Add1~18\,
	sumout => \TheRxFsk|Lowpass|Add1~21_sumout\,
	cout => \TheRxFsk|Lowpass|Add1~22\);

-- Location: LABCELL_X27_Y64_N33
\TheRxFsk|Lowpass|vNextWriteAddress~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|vNextWriteAddress~3_combout\ = ( \TheRxFsk|Lowpass|R.WriteAddress\(2) & ( \TheRxFsk|Lowpass|Add1~21_sumout\ ) ) # ( !\TheRxFsk|Lowpass|R.WriteAddress\(2) & ( (\TheRxFsk|Lowpass|Add1~21_sumout\ & (((!\TheRxFsk|Lowpass|R.WriteAddress\(1)) 
-- # (!\TheRxFsk|Lowpass|Equal2~0_combout\)) # (\TheRxFsk|Lowpass|R.WriteAddress\(0)))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001100110001001100110011000100110011001100110011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_R.WriteAddress\(0),
	datab => \TheRxFsk|Lowpass|ALT_INV_Add1~21_sumout\,
	datac => \TheRxFsk|Lowpass|ALT_INV_R.WriteAddress\(1),
	datad => \TheRxFsk|Lowpass|ALT_INV_Equal2~0_combout\,
	dataf => \TheRxFsk|Lowpass|ALT_INV_R.WriteAddress\(2),
	combout => \TheRxFsk|Lowpass|vNextWriteAddress~3_combout\);

-- Location: FF_X27_Y64_N34
\TheRxFsk|Lowpass|R.WriteAddress[5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|vNextWriteAddress~3_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	ena => \TheRxFsk|Lowpass|R.WriteAddress[0]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|R.WriteAddress\(5));

-- Location: LABCELL_X27_Y64_N18
\TheRxFsk|Lowpass|Add1~25\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add1~25_sumout\ = SUM(( !\TheRxFsk|Lowpass|R.WriteAddress\(6) ) + ( VCC ) + ( \TheRxFsk|Lowpass|Add1~22\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000000000001111000011110000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Lowpass|ALT_INV_R.WriteAddress\(6),
	cin => \TheRxFsk|Lowpass|Add1~22\,
	sumout => \TheRxFsk|Lowpass|Add1~25_sumout\);

-- Location: LABCELL_X27_Y64_N30
\TheRxFsk|Lowpass|R.WriteAddress[6]~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|R.WriteAddress[6]~3_combout\ = ( !\TheRxFsk|Lowpass|Add1~25_sumout\ )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111111111111111111111111111100000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \TheRxFsk|Lowpass|ALT_INV_Add1~25_sumout\,
	combout => \TheRxFsk|Lowpass|R.WriteAddress[6]~3_combout\);

-- Location: FF_X27_Y64_N31
\TheRxFsk|Lowpass|R.WriteAddress[6]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|R.WriteAddress[6]~3_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	ena => \TheRxFsk|Lowpass|R.WriteAddress[0]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|R.WriteAddress\(6));

-- Location: LABCELL_X27_Y64_N36
\TheRxFsk|Lowpass|Equal2~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Equal2~0_combout\ = ( !\TheRxFsk|Lowpass|R.WriteAddress\(4) & ( (!\TheRxFsk|Lowpass|R.WriteAddress\(5) & (\TheRxFsk|Lowpass|R.WriteAddress\(6) & \TheRxFsk|Lowpass|R.WriteAddress\(3))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000001100000000000000110000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Lowpass|ALT_INV_R.WriteAddress\(5),
	datac => \TheRxFsk|Lowpass|ALT_INV_R.WriteAddress\(6),
	datad => \TheRxFsk|Lowpass|ALT_INV_R.WriteAddress\(3),
	dataf => \TheRxFsk|Lowpass|ALT_INV_R.WriteAddress\(4),
	combout => \TheRxFsk|Lowpass|Equal2~0_combout\);

-- Location: LABCELL_X27_Y64_N24
\TheRxFsk|Lowpass|vNextWriteAddress~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|vNextWriteAddress~0_combout\ = ( \TheRxFsk|Lowpass|R.WriteAddress\(2) & ( !\TheRxFsk|Lowpass|R.WriteAddress\(0) ) ) # ( !\TheRxFsk|Lowpass|R.WriteAddress\(2) & ( (!\TheRxFsk|Lowpass|R.WriteAddress\(0) & 
-- ((!\TheRxFsk|Lowpass|R.WriteAddress\(1)) # (!\TheRxFsk|Lowpass|Equal2~0_combout\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111110000000000111111000000000011111111000000001111111100000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Lowpass|ALT_INV_R.WriteAddress\(1),
	datac => \TheRxFsk|Lowpass|ALT_INV_Equal2~0_combout\,
	datad => \TheRxFsk|Lowpass|ALT_INV_R.WriteAddress\(0),
	dataf => \TheRxFsk|Lowpass|ALT_INV_R.WriteAddress\(2),
	combout => \TheRxFsk|Lowpass|vNextWriteAddress~0_combout\);

-- Location: FF_X27_Y64_N25
\TheRxFsk|Lowpass|R.WriteAddress[0]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|vNextWriteAddress~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	ena => \TheRxFsk|Lowpass|R.WriteAddress[0]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|R.WriteAddress[0]~DUPLICATE_q\);

-- Location: FF_X27_Y64_N43
\TheRxFsk|Lowpass|R.WriteAddress[1]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|R.WriteAddress[1]~1_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	ena => \TheRxFsk|Lowpass|R.WriteAddress[0]~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|R.WriteAddress[1]~DUPLICATE_q\);

-- Location: MLABCELL_X25_Y64_N21
\TheRxFsk|Lowpass|R.WriteAddress[1]~_wirecell\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|R.WriteAddress[1]~_wirecell_combout\ = !\TheRxFsk|Lowpass|R.WriteAddress[1]~DUPLICATE_q\

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111000011110000111100001111000011110000111100001111000011110000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Lowpass|ALT_INV_R.WriteAddress[1]~DUPLICATE_q\,
	combout => \TheRxFsk|Lowpass|R.WriteAddress[1]~_wirecell_combout\);

-- Location: LABCELL_X27_Y64_N57
\TheRxFsk|Lowpass|R.WriteAddress[3]~_wirecell\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|R.WriteAddress[3]~_wirecell_combout\ = !\TheRxFsk|Lowpass|R.WriteAddress\(3)

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111100000000111111110000000011111111000000001111111100000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \TheRxFsk|Lowpass|ALT_INV_R.WriteAddress\(3),
	combout => \TheRxFsk|Lowpass|R.WriteAddress[3]~_wirecell_combout\);

-- Location: MLABCELL_X25_Y64_N0
\TheRxFsk|Lowpass|R.WriteAddress[6]~_wirecell\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|R.WriteAddress[6]~_wirecell_combout\ = ( !\TheRxFsk|Lowpass|R.WriteAddress\(6) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111111111111111111111111111100000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \TheRxFsk|Lowpass|ALT_INV_R.WriteAddress\(6),
	combout => \TheRxFsk|Lowpass|R.WriteAddress[6]~_wirecell_combout\);

-- Location: MLABCELL_X28_Y64_N0
\TheRxFsk|Lowpass|Add0~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add0~2\ = CARRY(( \TheRxFsk|Lowpass|R.ReadAddressSample[0]~DUPLICATE_q\ ) + ( VCC ) + ( !VCC ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressSample[0]~DUPLICATE_q\,
	cin => GND,
	cout => \TheRxFsk|Lowpass|Add0~2\);

-- Location: MLABCELL_X28_Y64_N3
\TheRxFsk|Lowpass|Add0~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add0~5_sumout\ = SUM(( \TheRxFsk|Lowpass|R.ReadAddressSample\(1) ) + ( GND ) + ( \TheRxFsk|Lowpass|Add0~2\ ))
-- \TheRxFsk|Lowpass|Add0~6\ = CARRY(( \TheRxFsk|Lowpass|R.ReadAddressSample\(1) ) + ( GND ) + ( \TheRxFsk|Lowpass|Add0~2\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000101010101010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressSample\(1),
	cin => \TheRxFsk|Lowpass|Add0~2\,
	sumout => \TheRxFsk|Lowpass|Add0~5_sumout\,
	cout => \TheRxFsk|Lowpass|Add0~6\);

-- Location: MLABCELL_X28_Y64_N6
\TheRxFsk|Lowpass|Add0~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add0~9_sumout\ = SUM(( \TheRxFsk|Lowpass|R.ReadAddressSample\(2) ) + ( GND ) + ( \TheRxFsk|Lowpass|Add0~6\ ))
-- \TheRxFsk|Lowpass|Add0~10\ = CARRY(( \TheRxFsk|Lowpass|R.ReadAddressSample\(2) ) + ( GND ) + ( \TheRxFsk|Lowpass|Add0~6\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressSample\(2),
	cin => \TheRxFsk|Lowpass|Add0~6\,
	sumout => \TheRxFsk|Lowpass|Add0~9_sumout\,
	cout => \TheRxFsk|Lowpass|Add0~10\);

-- Location: FF_X28_Y64_N8
\TheRxFsk|Lowpass|R.ReadAddressSample[2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|Add0~9_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	ena => \TheRxFsk|Lowpass|R.AddressState~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|R.ReadAddressSample\(2));

-- Location: FF_X28_Y64_N35
\TheRxFsk|Lowpass|R.ReadAddressSample[0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|NextR~6_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	ena => \TheRxFsk|Lowpass|R.AddressState~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|R.ReadAddressSample\(0));

-- Location: MLABCELL_X28_Y64_N9
\TheRxFsk|Lowpass|Add0~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add0~13_sumout\ = SUM(( \TheRxFsk|Lowpass|R.ReadAddressSample\(3) ) + ( GND ) + ( \TheRxFsk|Lowpass|Add0~10\ ))
-- \TheRxFsk|Lowpass|Add0~14\ = CARRY(( \TheRxFsk|Lowpass|R.ReadAddressSample\(3) ) + ( GND ) + ( \TheRxFsk|Lowpass|Add0~10\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressSample\(3),
	cin => \TheRxFsk|Lowpass|Add0~10\,
	sumout => \TheRxFsk|Lowpass|Add0~13_sumout\,
	cout => \TheRxFsk|Lowpass|Add0~14\);

-- Location: MLABCELL_X28_Y64_N54
\TheRxFsk|Lowpass|NextR~8\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|NextR~8_combout\ = ( \TheRxFsk|Lowpass|Equal0~0_combout\ & ( (\TheRxFsk|Lowpass|Add0~13_sumout\ & ((!\TheRxFsk|Lowpass|R.ReadAddressSample\(1)) # ((\TheRxFsk|Lowpass|R.ReadAddressSample\(0)) # 
-- (\TheRxFsk|Lowpass|R.ReadAddressSample\(2))))) ) ) # ( !\TheRxFsk|Lowpass|Equal0~0_combout\ & ( \TheRxFsk|Lowpass|Add0~13_sumout\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011111111000000001111111100000000101111110000000010111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressSample\(1),
	datab => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressSample\(2),
	datac => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressSample\(0),
	datad => \TheRxFsk|Lowpass|ALT_INV_Add0~13_sumout\,
	dataf => \TheRxFsk|Lowpass|ALT_INV_Equal0~0_combout\,
	combout => \TheRxFsk|Lowpass|NextR~8_combout\);

-- Location: FF_X28_Y64_N55
\TheRxFsk|Lowpass|R.ReadAddressSample[3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|NextR~8_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	ena => \TheRxFsk|Lowpass|R.AddressState~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|R.ReadAddressSample\(3));

-- Location: MLABCELL_X28_Y64_N12
\TheRxFsk|Lowpass|Add0~17\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add0~17_sumout\ = SUM(( \TheRxFsk|Lowpass|R.ReadAddressSample\(4) ) + ( GND ) + ( \TheRxFsk|Lowpass|Add0~14\ ))
-- \TheRxFsk|Lowpass|Add0~18\ = CARRY(( \TheRxFsk|Lowpass|R.ReadAddressSample\(4) ) + ( GND ) + ( \TheRxFsk|Lowpass|Add0~14\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressSample\(4),
	cin => \TheRxFsk|Lowpass|Add0~14\,
	sumout => \TheRxFsk|Lowpass|Add0~17_sumout\,
	cout => \TheRxFsk|Lowpass|Add0~18\);

-- Location: FF_X28_Y64_N13
\TheRxFsk|Lowpass|R.ReadAddressSample[4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|Add0~17_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	ena => \TheRxFsk|Lowpass|R.AddressState~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|R.ReadAddressSample\(4));

-- Location: MLABCELL_X28_Y64_N15
\TheRxFsk|Lowpass|Add0~21\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add0~21_sumout\ = SUM(( \TheRxFsk|Lowpass|R.ReadAddressSample\(5) ) + ( GND ) + ( \TheRxFsk|Lowpass|Add0~18\ ))
-- \TheRxFsk|Lowpass|Add0~22\ = CARRY(( \TheRxFsk|Lowpass|R.ReadAddressSample\(5) ) + ( GND ) + ( \TheRxFsk|Lowpass|Add0~18\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressSample\(5),
	cin => \TheRxFsk|Lowpass|Add0~18\,
	sumout => \TheRxFsk|Lowpass|Add0~21_sumout\,
	cout => \TheRxFsk|Lowpass|Add0~22\);

-- Location: FF_X28_Y64_N16
\TheRxFsk|Lowpass|R.ReadAddressSample[5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|Add0~21_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	ena => \TheRxFsk|Lowpass|R.AddressState~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|R.ReadAddressSample\(5));

-- Location: MLABCELL_X28_Y64_N18
\TheRxFsk|Lowpass|Add0~25\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add0~25_sumout\ = SUM(( \TheRxFsk|Lowpass|R.ReadAddressSample\(6) ) + ( GND ) + ( \TheRxFsk|Lowpass|Add0~22\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressSample\(6),
	cin => \TheRxFsk|Lowpass|Add0~22\,
	sumout => \TheRxFsk|Lowpass|Add0~25_sumout\);

-- Location: MLABCELL_X28_Y64_N57
\TheRxFsk|Lowpass|NextR~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|NextR~9_combout\ = ( \TheRxFsk|Lowpass|R.ReadAddressSample[0]~DUPLICATE_q\ & ( \TheRxFsk|Lowpass|Add0~25_sumout\ ) ) # ( !\TheRxFsk|Lowpass|R.ReadAddressSample[0]~DUPLICATE_q\ & ( (\TheRxFsk|Lowpass|Add0~25_sumout\ & 
-- ((!\TheRxFsk|Lowpass|R.ReadAddressSample\(1)) # ((!\TheRxFsk|Lowpass|Equal0~0_combout\) # (\TheRxFsk|Lowpass|R.ReadAddressSample\(2))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011111011000000001111101100000000111111110000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressSample\(1),
	datab => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressSample\(2),
	datac => \TheRxFsk|Lowpass|ALT_INV_Equal0~0_combout\,
	datad => \TheRxFsk|Lowpass|ALT_INV_Add0~25_sumout\,
	dataf => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressSample[0]~DUPLICATE_q\,
	combout => \TheRxFsk|Lowpass|NextR~9_combout\);

-- Location: FF_X28_Y64_N58
\TheRxFsk|Lowpass|R.ReadAddressSample[6]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|NextR~9_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	ena => \TheRxFsk|Lowpass|R.AddressState~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|R.ReadAddressSample\(6));

-- Location: MLABCELL_X28_Y64_N30
\TheRxFsk|Lowpass|Equal0~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Equal0~0_combout\ = ( !\TheRxFsk|Lowpass|R.ReadAddressSample\(4) & ( (\TheRxFsk|Lowpass|R.ReadAddressSample\(6) & (!\TheRxFsk|Lowpass|R.ReadAddressSample\(5) & \TheRxFsk|Lowpass|R.ReadAddressSample\(3))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000110000000000000011000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressSample\(6),
	datac => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressSample\(5),
	datad => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressSample\(3),
	dataf => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressSample\(4),
	combout => \TheRxFsk|Lowpass|Equal0~0_combout\);

-- Location: MLABCELL_X28_Y64_N24
\TheRxFsk|Lowpass|NextR~7\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|NextR~7_combout\ = ( \TheRxFsk|Lowpass|Equal0~0_combout\ & ( (\TheRxFsk|Lowpass|Add0~5_sumout\ & (((!\TheRxFsk|Lowpass|R.ReadAddressSample\(1)) # (\TheRxFsk|Lowpass|R.ReadAddressSample\(0))) # 
-- (\TheRxFsk|Lowpass|R.ReadAddressSample\(2)))) ) ) # ( !\TheRxFsk|Lowpass|Equal0~0_combout\ & ( \TheRxFsk|Lowpass|Add0~5_sumout\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010101010101010101010101010101010101000101010101010100010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_Add0~5_sumout\,
	datab => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressSample\(2),
	datac => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressSample\(0),
	datad => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressSample\(1),
	dataf => \TheRxFsk|Lowpass|ALT_INV_Equal0~0_combout\,
	combout => \TheRxFsk|Lowpass|NextR~7_combout\);

-- Location: FF_X28_Y64_N26
\TheRxFsk|Lowpass|R.ReadAddressSample[1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|NextR~7_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	ena => \TheRxFsk|Lowpass|R.AddressState~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|R.ReadAddressSample\(1));

-- Location: MLABCELL_X28_Y64_N33
\TheRxFsk|Lowpass|NextR~6\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|NextR~6_combout\ = ( \TheRxFsk|Lowpass|Equal0~0_combout\ & ( (!\TheRxFsk|Lowpass|R.ReadAddressSample\(0) & ((!\TheRxFsk|Lowpass|R.ReadAddressSample\(1)) # (\TheRxFsk|Lowpass|R.ReadAddressSample\(2)))) ) ) # ( 
-- !\TheRxFsk|Lowpass|Equal0~0_combout\ & ( !\TheRxFsk|Lowpass|R.ReadAddressSample\(0) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111100000000111111110000000010101111000000001010111100000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressSample\(1),
	datac => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressSample\(2),
	datad => \TheRxFsk|Lowpass|ALT_INV_R.ReadAddressSample\(0),
	dataf => \TheRxFsk|Lowpass|ALT_INV_Equal0~0_combout\,
	combout => \TheRxFsk|Lowpass|NextR~6_combout\);

-- Location: FF_X28_Y64_N34
\TheRxFsk|Lowpass|R.ReadAddressSample[0]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|NextR~6_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	ena => \TheRxFsk|Lowpass|R.AddressState~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|R.ReadAddressSample[0]~DUPLICATE_q\);

-- Location: FF_X28_Y64_N25
\TheRxFsk|Lowpass|R.ReadAddressSample[1]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|NextR~7_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	ena => \TheRxFsk|Lowpass|R.AddressState~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|R.ReadAddressSample[1]~DUPLICATE_q\);

-- Location: LABCELL_X17_Y64_N0
\TheRxFsk|Substracted[-14]~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Substracted[-14]~1_combout\ = ( \TheRxFsk|Add2~13_sumout\ & ( (!\TheRxFsk|Add2~5_sumout\) # (\TheRxFsk|Add2~1_sumout\) ) ) # ( !\TheRxFsk|Add2~13_sumout\ & ( (!\TheRxFsk|Add2~5_sumout\ & \TheRxFsk|Add2~1_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0010001000100010001000100010001010111011101110111011101110111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|ALT_INV_Add2~5_sumout\,
	datab => \TheRxFsk|ALT_INV_Add2~1_sumout\,
	dataf => \TheRxFsk|ALT_INV_Add2~13_sumout\,
	combout => \TheRxFsk|Substracted[-14]~1_combout\);

-- Location: LABCELL_X17_Y64_N3
\TheRxFsk|Substracted[-13]~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Substracted[-13]~2_combout\ = ( \TheRxFsk|Add2~17_sumout\ & ( (!\TheRxFsk|Add2~5_sumout\) # (\TheRxFsk|Add2~1_sumout\) ) ) # ( !\TheRxFsk|Add2~17_sumout\ & ( (!\TheRxFsk|Add2~5_sumout\ & \TheRxFsk|Add2~1_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0010001000100010001000100010001010111011101110111011101110111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|ALT_INV_Add2~5_sumout\,
	datab => \TheRxFsk|ALT_INV_Add2~1_sumout\,
	dataf => \TheRxFsk|ALT_INV_Add2~17_sumout\,
	combout => \TheRxFsk|Substracted[-13]~2_combout\);

-- Location: LABCELL_X17_Y64_N42
\TheRxFsk|Substracted[-12]~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Substracted[-12]~3_combout\ = ( \TheRxFsk|Add2~1_sumout\ & ( (!\TheRxFsk|Add2~5_sumout\) # (\TheRxFsk|Add2~21_sumout\) ) ) # ( !\TheRxFsk|Add2~1_sumout\ & ( (!\TheRxFsk|Add2~5_sumout\ & \TheRxFsk|Add2~21_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000101000001010000010100000101010101111101011111010111110101111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|ALT_INV_Add2~5_sumout\,
	datac => \TheRxFsk|ALT_INV_Add2~21_sumout\,
	dataf => \TheRxFsk|ALT_INV_Add2~1_sumout\,
	combout => \TheRxFsk|Substracted[-12]~3_combout\);

-- Location: LABCELL_X17_Y64_N45
\TheRxFsk|Substracted[-11]~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Substracted[-11]~4_combout\ = ( \TheRxFsk|Add2~25_sumout\ & ( (!\TheRxFsk|Add2~5_sumout\) # (\TheRxFsk|Add2~1_sumout\) ) ) # ( !\TheRxFsk|Add2~25_sumout\ & ( (!\TheRxFsk|Add2~5_sumout\ & \TheRxFsk|Add2~1_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0010001000100010001000100010001010111011101110111011101110111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|ALT_INV_Add2~5_sumout\,
	datab => \TheRxFsk|ALT_INV_Add2~1_sumout\,
	dataf => \TheRxFsk|ALT_INV_Add2~25_sumout\,
	combout => \TheRxFsk|Substracted[-11]~4_combout\);

-- Location: LABCELL_X17_Y64_N12
\TheRxFsk|Substracted[-10]~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Substracted[-10]~5_combout\ = ( \TheRxFsk|Add2~1_sumout\ & ( (!\TheRxFsk|Add2~5_sumout\) # (\TheRxFsk|Add2~29_sumout\) ) ) # ( !\TheRxFsk|Add2~1_sumout\ & ( (!\TheRxFsk|Add2~5_sumout\ & \TheRxFsk|Add2~29_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000101000001010000010100000101010101111101011111010111110101111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|ALT_INV_Add2~5_sumout\,
	datac => \TheRxFsk|ALT_INV_Add2~29_sumout\,
	dataf => \TheRxFsk|ALT_INV_Add2~1_sumout\,
	combout => \TheRxFsk|Substracted[-10]~5_combout\);

-- Location: LABCELL_X17_Y64_N15
\TheRxFsk|Substracted[-9]~6\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Substracted[-9]~6_combout\ = ( \TheRxFsk|Add2~1_sumout\ & ( (!\TheRxFsk|Add2~5_sumout\) # (\TheRxFsk|Add2~33_sumout\) ) ) # ( !\TheRxFsk|Add2~1_sumout\ & ( (!\TheRxFsk|Add2~5_sumout\ & \TheRxFsk|Add2~33_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000010101010000000001010101010101010111111111010101011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|ALT_INV_Add2~5_sumout\,
	datad => \TheRxFsk|ALT_INV_Add2~33_sumout\,
	dataf => \TheRxFsk|ALT_INV_Add2~1_sumout\,
	combout => \TheRxFsk|Substracted[-9]~6_combout\);

-- Location: LABCELL_X17_Y64_N30
\TheRxFsk|Substracted[-8]~7\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Substracted[-8]~7_combout\ = ( \TheRxFsk|Add2~37_sumout\ & ( (!\TheRxFsk|Add2~5_sumout\) # (\TheRxFsk|Add2~1_sumout\) ) ) # ( !\TheRxFsk|Add2~37_sumout\ & ( (!\TheRxFsk|Add2~5_sumout\ & \TheRxFsk|Add2~1_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0010001000100010001000100010001010111011101110111011101110111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|ALT_INV_Add2~5_sumout\,
	datab => \TheRxFsk|ALT_INV_Add2~1_sumout\,
	dataf => \TheRxFsk|ALT_INV_Add2~37_sumout\,
	combout => \TheRxFsk|Substracted[-8]~7_combout\);

-- Location: LABCELL_X17_Y64_N33
\TheRxFsk|Substracted[-7]~8\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Substracted[-7]~8_combout\ = ( \TheRxFsk|Add2~41_sumout\ & ( (!\TheRxFsk|Add2~5_sumout\) # (\TheRxFsk|Add2~1_sumout\) ) ) # ( !\TheRxFsk|Add2~41_sumout\ & ( (!\TheRxFsk|Add2~5_sumout\ & \TheRxFsk|Add2~1_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0010001000100010001000100010001010111011101110111011101110111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|ALT_INV_Add2~5_sumout\,
	datab => \TheRxFsk|ALT_INV_Add2~1_sumout\,
	dataf => \TheRxFsk|ALT_INV_Add2~41_sumout\,
	combout => \TheRxFsk|Substracted[-7]~8_combout\);

-- Location: LABCELL_X17_Y64_N48
\TheRxFsk|Substracted[-6]~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Substracted[-6]~9_combout\ = ( \TheRxFsk|Add2~45_sumout\ & ( (!\TheRxFsk|Add2~5_sumout\) # (\TheRxFsk|Add2~1_sumout\) ) ) # ( !\TheRxFsk|Add2~45_sumout\ & ( (!\TheRxFsk|Add2~5_sumout\ & \TheRxFsk|Add2~1_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0010001000100010001000100010001010111011101110111011101110111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|ALT_INV_Add2~5_sumout\,
	datab => \TheRxFsk|ALT_INV_Add2~1_sumout\,
	dataf => \TheRxFsk|ALT_INV_Add2~45_sumout\,
	combout => \TheRxFsk|Substracted[-6]~9_combout\);

-- Location: LABCELL_X17_Y64_N51
\TheRxFsk|Substracted[-5]~10\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Substracted[-5]~10_combout\ = ( \TheRxFsk|Add2~49_sumout\ & ( (!\TheRxFsk|Add2~5_sumout\) # (\TheRxFsk|Add2~1_sumout\) ) ) # ( !\TheRxFsk|Add2~49_sumout\ & ( (!\TheRxFsk|Add2~5_sumout\ & \TheRxFsk|Add2~1_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0010001000100010001000100010001010111011101110111011101110111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|ALT_INV_Add2~5_sumout\,
	datab => \TheRxFsk|ALT_INV_Add2~1_sumout\,
	dataf => \TheRxFsk|ALT_INV_Add2~49_sumout\,
	combout => \TheRxFsk|Substracted[-5]~10_combout\);

-- Location: LABCELL_X17_Y64_N54
\TheRxFsk|Substracted[-4]~11\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Substracted[-4]~11_combout\ = ( \TheRxFsk|Add2~53_sumout\ & ( (!\TheRxFsk|Add2~5_sumout\) # (\TheRxFsk|Add2~1_sumout\) ) ) # ( !\TheRxFsk|Add2~53_sumout\ & ( (!\TheRxFsk|Add2~5_sumout\ & \TheRxFsk|Add2~1_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0010001000100010001000100010001010111011101110111011101110111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|ALT_INV_Add2~5_sumout\,
	datab => \TheRxFsk|ALT_INV_Add2~1_sumout\,
	dataf => \TheRxFsk|ALT_INV_Add2~53_sumout\,
	combout => \TheRxFsk|Substracted[-4]~11_combout\);

-- Location: LABCELL_X17_Y64_N57
\TheRxFsk|Substracted[-3]~12\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Substracted[-3]~12_combout\ = (!\TheRxFsk|Add2~5_sumout\ & ((\TheRxFsk|Add2~57_sumout\) # (\TheRxFsk|Add2~1_sumout\))) # (\TheRxFsk|Add2~5_sumout\ & (\TheRxFsk|Add2~1_sumout\ & \TheRxFsk|Add2~57_sumout\))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0010101100101011001010110010101100101011001010110010101100101011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|ALT_INV_Add2~5_sumout\,
	datab => \TheRxFsk|ALT_INV_Add2~1_sumout\,
	datac => \TheRxFsk|ALT_INV_Add2~57_sumout\,
	combout => \TheRxFsk|Substracted[-3]~12_combout\);

-- Location: LABCELL_X17_Y64_N36
\TheRxFsk|Substracted[-2]~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Substracted[-2]~13_combout\ = ( \TheRxFsk|Add2~61_sumout\ & ( (!\TheRxFsk|Add2~5_sumout\) # (\TheRxFsk|Add2~1_sumout\) ) ) # ( !\TheRxFsk|Add2~61_sumout\ & ( (!\TheRxFsk|Add2~5_sumout\ & \TheRxFsk|Add2~1_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0010001000100010001000100010001010111011101110111011101110111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|ALT_INV_Add2~5_sumout\,
	datab => \TheRxFsk|ALT_INV_Add2~1_sumout\,
	dataf => \TheRxFsk|ALT_INV_Add2~61_sumout\,
	combout => \TheRxFsk|Substracted[-2]~13_combout\);

-- Location: LABCELL_X17_Y64_N39
\TheRxFsk|Substracted[-1]~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Substracted[-1]~14_combout\ = ( \TheRxFsk|Add2~65_sumout\ & ( (!\TheRxFsk|Add2~5_sumout\) # (\TheRxFsk|Add2~1_sumout\) ) ) # ( !\TheRxFsk|Add2~65_sumout\ & ( (!\TheRxFsk|Add2~5_sumout\ & \TheRxFsk|Add2~1_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0010001000100010001000100010001010111011101110111011101110111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|ALT_INV_Add2~5_sumout\,
	datab => \TheRxFsk|ALT_INV_Add2~1_sumout\,
	dataf => \TheRxFsk|ALT_INV_Add2~65_sumout\,
	combout => \TheRxFsk|Substracted[-1]~14_combout\);

-- Location: M10K_X26_Y64_N0
\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a0\ : cyclonev_ram_block
-- pragma translate_off
GENERIC MAP (
	mem_init2 => "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	mem_init1 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	mem_init0 => "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
	data_interleave_offset_in_bits => 1,
	data_interleave_width_in_bits => 1,
	init_file => "db/TbdRxFskBasic.ram0_DspFir_7e69c349.hdl.mif",
	init_file_layout => "port_a",
	logical_ram_name => "RxFsk:TheRxFsk|DspFir:Lowpass|altsyncram:SampleMemory_rtl_0|altsyncram_97s1:auto_generated|ALTSYNCRAM",
	mixed_port_feed_through_mode => "old",
	operation_mode => "dual_port",
	port_a_address_clear => "none",
	port_a_address_width => 7,
	port_a_byte_enable_clock => "none",
	port_a_data_out_clear => "none",
	port_a_data_out_clock => "none",
	port_a_data_width => 40,
	port_a_first_address => 0,
	port_a_first_bit_number => 0,
	port_a_last_address => 127,
	port_a_logical_ram_depth => 75,
	port_a_logical_ram_width => 16,
	port_a_read_during_write_mode => "new_data_no_nbe_read",
	port_b_address_clear => "none",
	port_b_address_clock => "clock0",
	port_b_address_width => 7,
	port_b_data_out_clear => "none",
	port_b_data_out_clock => "none",
	port_b_data_width => 40,
	port_b_first_address => 0,
	port_b_first_bit_number => 0,
	port_b_last_address => 127,
	port_b_logical_ram_depth => 75,
	port_b_logical_ram_width => 16,
	port_b_read_during_write_mode => "new_data_no_nbe_read",
	port_b_read_enable_clock => "clock0",
	ram_block_type => "M20K")
-- pragma translate_on
PORT MAP (
	portawe => \TheRxFsk|Bandpasses:11:Bandpass0|R.ValWet~q\,
	portbre => VCC,
	clk0 => \iClk~inputCLKENA0_outclk\,
	portadatain => \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTADATAIN_bus\,
	portaaddr => \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTAADDR_bus\,
	portbaddr => \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBADDR_bus\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	portbdataout => \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a0_PORTBDATAOUT_bus\);

-- Location: FF_X27_Y64_N41
\TheRxFsk|Lowpass|R.FirstSample\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	asdata => \TheRxFsk|Lowpass|R.AddressState~q\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|R.FirstSample~q\);

-- Location: LABCELL_X24_Y64_N57
\TheRxFsk|Add2~5_wirecell\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Add2~5_wirecell_combout\ = !\TheRxFsk|Add2~5_sumout\

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1010101010101010101010101010101010101010101010101010101010101010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|ALT_INV_Add2~5_sumout\,
	combout => \TheRxFsk|Add2~5_wirecell_combout\);

-- Location: LABCELL_X24_Y64_N54
\TheRxFsk|result~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|result~0_combout\ = ( \TheRxFsk|Add2~1_sumout\ & ( !\TheRxFsk|Add2~5_sumout\ ) ) # ( !\TheRxFsk|Add2~1_sumout\ & ( \TheRxFsk|Add2~5_sumout\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010101010101010101010101010110101010101010101010101010101010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|ALT_INV_Add2~5_sumout\,
	dataf => \TheRxFsk|ALT_INV_Add2~1_sumout\,
	combout => \TheRxFsk|result~0_combout\);

-- Location: FF_X24_Y64_N4
\TheRxFsk|Lowpass|DdryDelayed[-15]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Add2~9_sumout\,
	asdata => \TheRxFsk|Add2~5_wirecell_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => \TheRxFsk|result~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|DdryDelayed[-15]~q\);

-- Location: MLABCELL_X25_Y64_N18
\TheRxFsk|Lowpass|Sample[-15]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Sample[-15]~0_combout\ = ( \TheRxFsk|Lowpass|DdryDelayed[-15]~q\ & ( (!\TheRxFsk|Lowpass|R.FirstSample~q\) # (\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a0~portbdataout\) ) ) # ( !\TheRxFsk|Lowpass|DdryDelayed[-15]~q\ 
-- & ( (\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a0~portbdataout\ & \TheRxFsk|Lowpass|R.FirstSample~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000001111000000000000111111111111000011111111111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a0~portbdataout\,
	datad => \TheRxFsk|Lowpass|ALT_INV_R.FirstSample~q\,
	dataf => \TheRxFsk|Lowpass|ALT_INV_DdryDelayed[-15]~q\,
	combout => \TheRxFsk|Lowpass|Sample[-15]~0_combout\);

-- Location: FF_X24_Y64_N7
\TheRxFsk|Lowpass|DdryDelayed[-14]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Add2~13_sumout\,
	asdata => \TheRxFsk|Add2~5_wirecell_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => \TheRxFsk|result~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|DdryDelayed[-14]~q\);

-- Location: MLABCELL_X25_Y64_N39
\TheRxFsk|Lowpass|Sample[-14]~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Sample[-14]~1_combout\ = ( \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a1\ & ( (\TheRxFsk|Lowpass|DdryDelayed[-14]~q\) # (\TheRxFsk|Lowpass|R.FirstSample~q\) ) ) # ( 
-- !\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a1\ & ( (!\TheRxFsk|Lowpass|R.FirstSample~q\ & \TheRxFsk|Lowpass|DdryDelayed[-14]~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011110000000000001111000000001111111111110000111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Lowpass|ALT_INV_R.FirstSample~q\,
	datad => \TheRxFsk|Lowpass|ALT_INV_DdryDelayed[-14]~q\,
	dataf => \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a1\,
	combout => \TheRxFsk|Lowpass|Sample[-14]~1_combout\);

-- Location: FF_X24_Y64_N10
\TheRxFsk|Lowpass|DdryDelayed[-13]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Add2~17_sumout\,
	asdata => \TheRxFsk|Add2~5_wirecell_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => \TheRxFsk|result~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|DdryDelayed[-13]~q\);

-- Location: LABCELL_X27_Y64_N54
\TheRxFsk|Lowpass|Sample[-13]~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Sample[-13]~2_combout\ = ( \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a2\ & ( (\TheRxFsk|Lowpass|DdryDelayed[-13]~q\) # (\TheRxFsk|Lowpass|R.FirstSample~q\) ) ) # ( 
-- !\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a2\ & ( (!\TheRxFsk|Lowpass|R.FirstSample~q\ & \TheRxFsk|Lowpass|DdryDelayed[-13]~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000110000001100000011000000110000111111001111110011111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Lowpass|ALT_INV_R.FirstSample~q\,
	datac => \TheRxFsk|Lowpass|ALT_INV_DdryDelayed[-13]~q\,
	dataf => \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a2\,
	combout => \TheRxFsk|Lowpass|Sample[-13]~2_combout\);

-- Location: FF_X24_Y64_N13
\TheRxFsk|Lowpass|DdryDelayed[-12]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Add2~21_sumout\,
	asdata => \TheRxFsk|Add2~5_wirecell_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => \TheRxFsk|result~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|DdryDelayed[-12]~q\);

-- Location: MLABCELL_X25_Y64_N3
\TheRxFsk|Lowpass|Sample[-12]~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Sample[-12]~3_combout\ = (!\TheRxFsk|Lowpass|R.FirstSample~q\ & ((\TheRxFsk|Lowpass|DdryDelayed[-12]~q\))) # (\TheRxFsk|Lowpass|R.FirstSample~q\ & (\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a3\))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010111110101000001011111010100000101111101010000010111110101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a3\,
	datac => \TheRxFsk|Lowpass|ALT_INV_R.FirstSample~q\,
	datad => \TheRxFsk|Lowpass|ALT_INV_DdryDelayed[-12]~q\,
	combout => \TheRxFsk|Lowpass|Sample[-12]~3_combout\);

-- Location: FF_X24_Y64_N16
\TheRxFsk|Lowpass|DdryDelayed[-11]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Add2~25_sumout\,
	asdata => \TheRxFsk|Add2~5_wirecell_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => \TheRxFsk|result~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|DdryDelayed[-11]~q\);

-- Location: LABCELL_X29_Y64_N27
\TheRxFsk|Lowpass|Sample[-11]~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Sample[-11]~4_combout\ = ( \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a4\ & ( (\TheRxFsk|Lowpass|DdryDelayed[-11]~q\) # (\TheRxFsk|Lowpass|R.FirstSample~q\) ) ) # ( 
-- !\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a4\ & ( (!\TheRxFsk|Lowpass|R.FirstSample~q\ & \TheRxFsk|Lowpass|DdryDelayed[-11]~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011110000000000001111000000001111111111110000111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Lowpass|ALT_INV_R.FirstSample~q\,
	datad => \TheRxFsk|Lowpass|ALT_INV_DdryDelayed[-11]~q\,
	dataf => \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a4\,
	combout => \TheRxFsk|Lowpass|Sample[-11]~4_combout\);

-- Location: FF_X24_Y64_N19
\TheRxFsk|Lowpass|DdryDelayed[-10]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Add2~29_sumout\,
	asdata => \TheRxFsk|Add2~5_wirecell_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => \TheRxFsk|result~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|DdryDelayed[-10]~q\);

-- Location: MLABCELL_X25_Y64_N15
\TheRxFsk|Lowpass|Sample[-10]~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Sample[-10]~5_combout\ = ( \TheRxFsk|Lowpass|DdryDelayed[-10]~q\ & ( (!\TheRxFsk|Lowpass|R.FirstSample~q\) # (\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a5\) ) ) # ( !\TheRxFsk|Lowpass|DdryDelayed[-10]~q\ & ( 
-- (\TheRxFsk|Lowpass|R.FirstSample~q\ & \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a5\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000001111000000000000111111110000111111111111000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Lowpass|ALT_INV_R.FirstSample~q\,
	datad => \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a5\,
	dataf => \TheRxFsk|Lowpass|ALT_INV_DdryDelayed[-10]~q\,
	combout => \TheRxFsk|Lowpass|Sample[-10]~5_combout\);

-- Location: FF_X24_Y64_N22
\TheRxFsk|Lowpass|DdryDelayed[-9]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Add2~33_sumout\,
	asdata => \TheRxFsk|Add2~5_wirecell_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => \TheRxFsk|result~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|DdryDelayed[-9]~q\);

-- Location: LABCELL_X29_Y64_N57
\TheRxFsk|Lowpass|Sample[-9]~6\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Sample[-9]~6_combout\ = ( \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a6\ & ( (\TheRxFsk|Lowpass|DdryDelayed[-9]~q\) # (\TheRxFsk|Lowpass|R.FirstSample~q\) ) ) # ( 
-- !\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a6\ & ( (!\TheRxFsk|Lowpass|R.FirstSample~q\ & \TheRxFsk|Lowpass|DdryDelayed[-9]~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011110000000000001111000000001111111111110000111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Lowpass|ALT_INV_R.FirstSample~q\,
	datad => \TheRxFsk|Lowpass|ALT_INV_DdryDelayed[-9]~q\,
	dataf => \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a6\,
	combout => \TheRxFsk|Lowpass|Sample[-9]~6_combout\);

-- Location: FF_X24_Y64_N25
\TheRxFsk|Lowpass|DdryDelayed[-8]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Add2~37_sumout\,
	asdata => \TheRxFsk|Add2~5_wirecell_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => \TheRxFsk|result~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|DdryDelayed[-8]~q\);

-- Location: LABCELL_X30_Y64_N36
\TheRxFsk|Lowpass|Sample[-8]~7\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Sample[-8]~7_combout\ = ( \TheRxFsk|Lowpass|R.FirstSample~q\ & ( \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a7\ ) ) # ( !\TheRxFsk|Lowpass|R.FirstSample~q\ & ( 
-- \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a7\ & ( \TheRxFsk|Lowpass|DdryDelayed[-8]~q\ ) ) ) # ( !\TheRxFsk|Lowpass|R.FirstSample~q\ & ( !\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a7\ & ( 
-- \TheRxFsk|Lowpass|DdryDelayed[-8]~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001100110011000000000000000000110011001100111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Lowpass|ALT_INV_DdryDelayed[-8]~q\,
	datae => \TheRxFsk|Lowpass|ALT_INV_R.FirstSample~q\,
	dataf => \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a7\,
	combout => \TheRxFsk|Lowpass|Sample[-8]~7_combout\);

-- Location: FF_X24_Y64_N28
\TheRxFsk|Lowpass|DdryDelayed[-7]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Add2~41_sumout\,
	asdata => \TheRxFsk|Add2~5_wirecell_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => \TheRxFsk|result~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|DdryDelayed[-7]~q\);

-- Location: MLABCELL_X25_Y64_N30
\TheRxFsk|Lowpass|Sample[-7]~8\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Sample[-7]~8_combout\ = (!\TheRxFsk|Lowpass|R.FirstSample~q\ & (\TheRxFsk|Lowpass|DdryDelayed[-7]~q\)) # (\TheRxFsk|Lowpass|R.FirstSample~q\ & ((\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a8\)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000110000111111000011000011111100001100001111110000110000111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Lowpass|ALT_INV_R.FirstSample~q\,
	datac => \TheRxFsk|Lowpass|ALT_INV_DdryDelayed[-7]~q\,
	datad => \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a8\,
	combout => \TheRxFsk|Lowpass|Sample[-7]~8_combout\);

-- Location: FF_X24_Y64_N31
\TheRxFsk|Lowpass|DdryDelayed[-6]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Add2~45_sumout\,
	asdata => \TheRxFsk|Add2~5_wirecell_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => \TheRxFsk|result~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|DdryDelayed[-6]~q\);

-- Location: MLABCELL_X25_Y64_N33
\TheRxFsk|Lowpass|Sample[-6]~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Sample[-6]~9_combout\ = ( \TheRxFsk|Lowpass|DdryDelayed[-6]~q\ & ( (!\TheRxFsk|Lowpass|R.FirstSample~q\) # (\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a9\) ) ) # ( !\TheRxFsk|Lowpass|DdryDelayed[-6]~q\ & ( 
-- (\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a9\ & \TheRxFsk|Lowpass|R.FirstSample~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000100010001000100010001000111011101110111011101110111011101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a9\,
	datab => \TheRxFsk|Lowpass|ALT_INV_R.FirstSample~q\,
	dataf => \TheRxFsk|Lowpass|ALT_INV_DdryDelayed[-6]~q\,
	combout => \TheRxFsk|Lowpass|Sample[-6]~9_combout\);

-- Location: FF_X24_Y64_N34
\TheRxFsk|Lowpass|DdryDelayed[-5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Add2~49_sumout\,
	asdata => \TheRxFsk|Add2~5_wirecell_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => \TheRxFsk|result~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|DdryDelayed[-5]~q\);

-- Location: MLABCELL_X25_Y64_N42
\TheRxFsk|Lowpass|Sample[-5]~10\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Sample[-5]~10_combout\ = ( \TheRxFsk|Lowpass|R.FirstSample~q\ & ( \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a10\ ) ) # ( !\TheRxFsk|Lowpass|R.FirstSample~q\ & ( 
-- \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a10\ & ( \TheRxFsk|Lowpass|DdryDelayed[-5]~q\ ) ) ) # ( !\TheRxFsk|Lowpass|R.FirstSample~q\ & ( !\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a10\ & ( 
-- \TheRxFsk|Lowpass|DdryDelayed[-5]~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001100110011000000000000000000110011001100111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Lowpass|ALT_INV_DdryDelayed[-5]~q\,
	datae => \TheRxFsk|Lowpass|ALT_INV_R.FirstSample~q\,
	dataf => \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a10\,
	combout => \TheRxFsk|Lowpass|Sample[-5]~10_combout\);

-- Location: FF_X24_Y64_N37
\TheRxFsk|Lowpass|DdryDelayed[-4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Add2~53_sumout\,
	asdata => \TheRxFsk|Add2~5_wirecell_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => \TheRxFsk|result~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|DdryDelayed[-4]~q\);

-- Location: MLABCELL_X25_Y64_N24
\TheRxFsk|Lowpass|Sample[-4]~11\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Sample[-4]~11_combout\ = ( \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a11\ & ( (\TheRxFsk|Lowpass|R.FirstSample~q\) # (\TheRxFsk|Lowpass|DdryDelayed[-4]~q\) ) ) # ( 
-- !\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a11\ & ( (\TheRxFsk|Lowpass|DdryDelayed[-4]~q\ & !\TheRxFsk|Lowpass|R.FirstSample~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100000000000011110000000000001111111111110000111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Lowpass|ALT_INV_DdryDelayed[-4]~q\,
	datad => \TheRxFsk|Lowpass|ALT_INV_R.FirstSample~q\,
	dataf => \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a11\,
	combout => \TheRxFsk|Lowpass|Sample[-4]~11_combout\);

-- Location: FF_X24_Y64_N40
\TheRxFsk|Lowpass|DdryDelayed[-3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Add2~57_sumout\,
	asdata => \TheRxFsk|Add2~5_wirecell_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => \TheRxFsk|result~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|DdryDelayed[-3]~q\);

-- Location: MLABCELL_X25_Y64_N54
\TheRxFsk|Lowpass|Sample[-3]~12\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Sample[-3]~12_combout\ = ( \TheRxFsk|Lowpass|DdryDelayed[-3]~q\ & ( (!\TheRxFsk|Lowpass|R.FirstSample~q\) # (\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a12\) ) ) # ( !\TheRxFsk|Lowpass|DdryDelayed[-3]~q\ & ( 
-- (\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a12\ & \TheRxFsk|Lowpass|R.FirstSample~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000110011000000000011001111111111001100111111111100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a12\,
	datad => \TheRxFsk|Lowpass|ALT_INV_R.FirstSample~q\,
	dataf => \TheRxFsk|Lowpass|ALT_INV_DdryDelayed[-3]~q\,
	combout => \TheRxFsk|Lowpass|Sample[-3]~12_combout\);

-- Location: FF_X24_Y64_N43
\TheRxFsk|Lowpass|DdryDelayed[-2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Add2~61_sumout\,
	asdata => \TheRxFsk|Add2~5_wirecell_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => \TheRxFsk|result~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|DdryDelayed[-2]~q\);

-- Location: LABCELL_X29_Y64_N12
\TheRxFsk|Lowpass|Sample[-2]~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Sample[-2]~13_combout\ = ( \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a13\ & ( (\TheRxFsk|Lowpass|DdryDelayed[-2]~q\) # (\TheRxFsk|Lowpass|R.FirstSample~q\) ) ) # ( 
-- !\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a13\ & ( (!\TheRxFsk|Lowpass|R.FirstSample~q\ & \TheRxFsk|Lowpass|DdryDelayed[-2]~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000110000001100000011000000110000111111001111110011111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Lowpass|ALT_INV_R.FirstSample~q\,
	datac => \TheRxFsk|Lowpass|ALT_INV_DdryDelayed[-2]~q\,
	dataf => \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a13\,
	combout => \TheRxFsk|Lowpass|Sample[-2]~13_combout\);

-- Location: FF_X24_Y64_N47
\TheRxFsk|Lowpass|DdryDelayed[-1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Add2~65_sumout\,
	asdata => \TheRxFsk|Add2~5_wirecell_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => \TheRxFsk|result~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|DdryDelayed[-1]~q\);

-- Location: LABCELL_X27_Y64_N27
\TheRxFsk|Lowpass|Sample[-1]~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Sample[-1]~14_combout\ = ( \TheRxFsk|Lowpass|R.FirstSample~q\ & ( \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a14\ ) ) # ( !\TheRxFsk|Lowpass|R.FirstSample~q\ & ( \TheRxFsk|Lowpass|DdryDelayed[-1]~q\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111000011110000111100000000111111110000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Lowpass|ALT_INV_DdryDelayed[-1]~q\,
	datad => \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a14\,
	dataf => \TheRxFsk|Lowpass|ALT_INV_R.FirstSample~q\,
	combout => \TheRxFsk|Lowpass|Sample[-1]~14_combout\);

-- Location: FF_X24_Y64_N49
\TheRxFsk|Lowpass|DdryDelayed[0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Add2~1_sumout\,
	asdata => \TheRxFsk|Add2~5_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => \TheRxFsk|result~0_combout\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|DdryDelayed\(0));

-- Location: LABCELL_X27_Y64_N39
\TheRxFsk|Lowpass|Sample[0]~15\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Sample[0]~15_combout\ = ( \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a15\ & ( (\TheRxFsk|Lowpass|R.FirstSample~q\) # (\TheRxFsk|Lowpass|DdryDelayed\(0)) ) ) # ( 
-- !\TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ram_block1a15\ & ( (\TheRxFsk|Lowpass|DdryDelayed\(0) & !\TheRxFsk|Lowpass|R.FirstSample~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100000000000011110000000000001111111111110000111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Lowpass|ALT_INV_DdryDelayed\(0),
	datad => \TheRxFsk|Lowpass|ALT_INV_R.FirstSample~q\,
	dataf => \TheRxFsk|Lowpass|SampleMemory_rtl_0|auto_generated|ALT_INV_ram_block1a15\,
	combout => \TheRxFsk|Lowpass|Sample[0]~15_combout\);

-- Location: DSP_X32_Y65_N0
\TheRxFsk|Lowpass|Mult0~8\ : cyclonev_mac
-- pragma translate_off
GENERIC MAP (
	accumulate_clock => "none",
	ax_clock => "0",
	ax_width => 18,
	ay_scan_in_clock => "none",
	ay_scan_in_width => 19,
	ay_use_scan_in => "false",
	az_clock => "none",
	bx_clock => "none",
	by_clock => "none",
	by_use_scan_in => "false",
	bz_clock => "none",
	coef_a_0 => 0,
	coef_a_1 => 0,
	coef_a_2 => 0,
	coef_a_3 => 0,
	coef_a_4 => 0,
	coef_a_5 => 0,
	coef_a_6 => 0,
	coef_a_7 => 0,
	coef_b_0 => 0,
	coef_b_1 => 0,
	coef_b_2 => 0,
	coef_b_3 => 0,
	coef_b_4 => 0,
	coef_b_5 => 0,
	coef_b_6 => 0,
	coef_b_7 => 0,
	coef_sel_a_clock => "none",
	coef_sel_b_clock => "none",
	delay_scan_out_ay => "false",
	delay_scan_out_by => "false",
	enable_double_accum => "false",
	load_const_clock => "none",
	load_const_value => 0,
	mode_sub_location => 0,
	negate_clock => "none",
	operand_source_max => "input",
	operand_source_may => "input",
	operand_source_mbx => "input",
	operand_source_mby => "input",
	operation_mode => "m18x18_full",
	output_clock => "none",
	preadder_subtract_a => "false",
	preadder_subtract_b => "false",
	result_a_width => 64,
	signed_max => "true",
	signed_may => "true",
	signed_mbx => "false",
	signed_mby => "false",
	sub_clock => "none",
	use_chainadder => "false")
-- pragma translate_on
PORT MAP (
	sub => GND,
	negate => GND,
	aclr => \TheRxFsk|Lowpass|Mult0~8_ACLR_bus\,
	clk => \TheRxFsk|Lowpass|Mult0~8_CLK_bus\,
	ena => \TheRxFsk|Lowpass|Mult0~8_ENA_bus\,
	ax => \TheRxFsk|Lowpass|Mult0~8_AX_bus\,
	ay => \TheRxFsk|Lowpass|Mult0~8_AY_bus\,
	resulta => \TheRxFsk|Lowpass|Mult0~8_RESULTA_bus\);

-- Location: LABCELL_X31_Y65_N48
\TheRxFsk|Lowpass|vAdd~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|vAdd~1_combout\ = ( !\TheRxFsk|Lowpass|Mult0~18\ & ( !\TheRxFsk|Lowpass|Mult0~14\ & ( (!\TheRxFsk|Lowpass|Mult0~17\ & (!\TheRxFsk|Lowpass|Mult0~9\ & (!\TheRxFsk|Lowpass|Mult0~15\ & !\TheRxFsk|Lowpass|Mult0~16\))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1000000000000000000000000000000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_Mult0~17\,
	datab => \TheRxFsk|Lowpass|ALT_INV_Mult0~9\,
	datac => \TheRxFsk|Lowpass|ALT_INV_Mult0~15\,
	datad => \TheRxFsk|Lowpass|ALT_INV_Mult0~16\,
	datae => \TheRxFsk|Lowpass|ALT_INV_Mult0~18\,
	dataf => \TheRxFsk|Lowpass|ALT_INV_Mult0~14\,
	combout => \TheRxFsk|Lowpass|vAdd~1_combout\);

-- Location: LABCELL_X31_Y65_N57
\TheRxFsk|Lowpass|vAdd~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|vAdd~2_combout\ = ( !\TheRxFsk|Lowpass|Mult0~11\ & ( !\TheRxFsk|Lowpass|Mult0~12\ & ( (!\TheRxFsk|Lowpass|Mult0~8_resulta\ & (!\TheRxFsk|Lowpass|Mult0~21\ & !\TheRxFsk|Lowpass|Mult0~10\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1010000000000000000000000000000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_Mult0~8_resulta\,
	datac => \TheRxFsk|Lowpass|ALT_INV_Mult0~21\,
	datad => \TheRxFsk|Lowpass|ALT_INV_Mult0~10\,
	datae => \TheRxFsk|Lowpass|ALT_INV_Mult0~11\,
	dataf => \TheRxFsk|Lowpass|ALT_INV_Mult0~12\,
	combout => \TheRxFsk|Lowpass|vAdd~2_combout\);

-- Location: LABCELL_X33_Y65_N54
\TheRxFsk|Lowpass|vAdd~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|vAdd~0_combout\ = ( \TheRxFsk|Lowpass|Mult0~20\ & ( \TheRxFsk|Lowpass|Mult0~13\ ) ) # ( !\TheRxFsk|Lowpass|Mult0~20\ & ( \TheRxFsk|Lowpass|Mult0~13\ ) ) # ( \TheRxFsk|Lowpass|Mult0~20\ & ( !\TheRxFsk|Lowpass|Mult0~13\ ) ) # ( 
-- !\TheRxFsk|Lowpass|Mult0~20\ & ( !\TheRxFsk|Lowpass|Mult0~13\ & ( ((!\TheRxFsk|Lowpass|vAdd~1_combout\) # ((!\TheRxFsk|Lowpass|vAdd~2_combout\) # (\TheRxFsk|Lowpass|Mult0~22\))) # (\TheRxFsk|Lowpass|Mult0~19\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111110111111111111111111111111111111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_Mult0~19\,
	datab => \TheRxFsk|Lowpass|ALT_INV_vAdd~1_combout\,
	datac => \TheRxFsk|Lowpass|ALT_INV_vAdd~2_combout\,
	datad => \TheRxFsk|Lowpass|ALT_INV_Mult0~22\,
	datae => \TheRxFsk|Lowpass|ALT_INV_Mult0~20\,
	dataf => \TheRxFsk|Lowpass|ALT_INV_Mult0~13\,
	combout => \TheRxFsk|Lowpass|vAdd~0_combout\);

-- Location: LABCELL_X33_Y65_N0
\TheRxFsk|Lowpass|Add3~69\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add3~69_sumout\ = SUM(( (\TheRxFsk|Lowpass|Mult0~39\ & \TheRxFsk|Lowpass|vAdd~0_combout\) ) + ( \TheRxFsk|Lowpass|Mult0~23\ ) + ( !VCC ))
-- \TheRxFsk|Lowpass|Add3~70\ = CARRY(( (\TheRxFsk|Lowpass|Mult0~39\ & \TheRxFsk|Lowpass|vAdd~0_combout\) ) + ( \TheRxFsk|Lowpass|Mult0~23\ ) + ( !VCC ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000001010101",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_Mult0~39\,
	datac => \TheRxFsk|Lowpass|ALT_INV_Mult0~23\,
	datad => \TheRxFsk|Lowpass|ALT_INV_vAdd~0_combout\,
	cin => GND,
	sumout => \TheRxFsk|Lowpass|Add3~69_sumout\,
	cout => \TheRxFsk|Lowpass|Add3~70\);

-- Location: LABCELL_X33_Y65_N3
\TheRxFsk|Lowpass|Add3~65\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add3~65_sumout\ = SUM(( GND ) + ( \TheRxFsk|Lowpass|Mult0~24\ ) + ( \TheRxFsk|Lowpass|Add3~70\ ))
-- \TheRxFsk|Lowpass|Add3~66\ = CARRY(( GND ) + ( \TheRxFsk|Lowpass|Mult0~24\ ) + ( \TheRxFsk|Lowpass|Add3~70\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Lowpass|ALT_INV_Mult0~24\,
	cin => \TheRxFsk|Lowpass|Add3~70\,
	sumout => \TheRxFsk|Lowpass|Add3~65_sumout\,
	cout => \TheRxFsk|Lowpass|Add3~66\);

-- Location: LABCELL_X33_Y65_N6
\TheRxFsk|Lowpass|Add3~61\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add3~61_sumout\ = SUM(( GND ) + ( \TheRxFsk|Lowpass|Mult0~25\ ) + ( \TheRxFsk|Lowpass|Add3~66\ ))
-- \TheRxFsk|Lowpass|Add3~62\ = CARRY(( GND ) + ( \TheRxFsk|Lowpass|Mult0~25\ ) + ( \TheRxFsk|Lowpass|Add3~66\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Lowpass|ALT_INV_Mult0~25\,
	cin => \TheRxFsk|Lowpass|Add3~66\,
	sumout => \TheRxFsk|Lowpass|Add3~61_sumout\,
	cout => \TheRxFsk|Lowpass|Add3~62\);

-- Location: LABCELL_X33_Y65_N9
\TheRxFsk|Lowpass|Add3~57\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add3~57_sumout\ = SUM(( GND ) + ( \TheRxFsk|Lowpass|Mult0~26\ ) + ( \TheRxFsk|Lowpass|Add3~62\ ))
-- \TheRxFsk|Lowpass|Add3~58\ = CARRY(( GND ) + ( \TheRxFsk|Lowpass|Mult0~26\ ) + ( \TheRxFsk|Lowpass|Add3~62\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Lowpass|ALT_INV_Mult0~26\,
	cin => \TheRxFsk|Lowpass|Add3~62\,
	sumout => \TheRxFsk|Lowpass|Add3~57_sumout\,
	cout => \TheRxFsk|Lowpass|Add3~58\);

-- Location: LABCELL_X33_Y65_N12
\TheRxFsk|Lowpass|Add3~53\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add3~53_sumout\ = SUM(( GND ) + ( \TheRxFsk|Lowpass|Mult0~27\ ) + ( \TheRxFsk|Lowpass|Add3~58\ ))
-- \TheRxFsk|Lowpass|Add3~54\ = CARRY(( GND ) + ( \TheRxFsk|Lowpass|Mult0~27\ ) + ( \TheRxFsk|Lowpass|Add3~58\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Lowpass|ALT_INV_Mult0~27\,
	cin => \TheRxFsk|Lowpass|Add3~58\,
	sumout => \TheRxFsk|Lowpass|Add3~53_sumout\,
	cout => \TheRxFsk|Lowpass|Add3~54\);

-- Location: LABCELL_X33_Y65_N15
\TheRxFsk|Lowpass|Add3~49\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add3~49_sumout\ = SUM(( \TheRxFsk|Lowpass|Mult0~28\ ) + ( GND ) + ( \TheRxFsk|Lowpass|Add3~54\ ))
-- \TheRxFsk|Lowpass|Add3~50\ = CARRY(( \TheRxFsk|Lowpass|Mult0~28\ ) + ( GND ) + ( \TheRxFsk|Lowpass|Add3~54\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \TheRxFsk|Lowpass|ALT_INV_Mult0~28\,
	cin => \TheRxFsk|Lowpass|Add3~54\,
	sumout => \TheRxFsk|Lowpass|Add3~49_sumout\,
	cout => \TheRxFsk|Lowpass|Add3~50\);

-- Location: LABCELL_X33_Y65_N18
\TheRxFsk|Lowpass|Add3~45\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add3~45_sumout\ = SUM(( GND ) + ( \TheRxFsk|Lowpass|Mult0~29\ ) + ( \TheRxFsk|Lowpass|Add3~50\ ))
-- \TheRxFsk|Lowpass|Add3~46\ = CARRY(( GND ) + ( \TheRxFsk|Lowpass|Mult0~29\ ) + ( \TheRxFsk|Lowpass|Add3~50\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Lowpass|ALT_INV_Mult0~29\,
	cin => \TheRxFsk|Lowpass|Add3~50\,
	sumout => \TheRxFsk|Lowpass|Add3~45_sumout\,
	cout => \TheRxFsk|Lowpass|Add3~46\);

-- Location: LABCELL_X33_Y65_N21
\TheRxFsk|Lowpass|Add3~41\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add3~41_sumout\ = SUM(( GND ) + ( \TheRxFsk|Lowpass|Mult0~30\ ) + ( \TheRxFsk|Lowpass|Add3~46\ ))
-- \TheRxFsk|Lowpass|Add3~42\ = CARRY(( GND ) + ( \TheRxFsk|Lowpass|Mult0~30\ ) + ( \TheRxFsk|Lowpass|Add3~46\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Lowpass|ALT_INV_Mult0~30\,
	cin => \TheRxFsk|Lowpass|Add3~46\,
	sumout => \TheRxFsk|Lowpass|Add3~41_sumout\,
	cout => \TheRxFsk|Lowpass|Add3~42\);

-- Location: LABCELL_X33_Y65_N24
\TheRxFsk|Lowpass|Add3~37\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add3~37_sumout\ = SUM(( GND ) + ( \TheRxFsk|Lowpass|Mult0~31\ ) + ( \TheRxFsk|Lowpass|Add3~42\ ))
-- \TheRxFsk|Lowpass|Add3~38\ = CARRY(( GND ) + ( \TheRxFsk|Lowpass|Mult0~31\ ) + ( \TheRxFsk|Lowpass|Add3~42\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Lowpass|ALT_INV_Mult0~31\,
	cin => \TheRxFsk|Lowpass|Add3~42\,
	sumout => \TheRxFsk|Lowpass|Add3~37_sumout\,
	cout => \TheRxFsk|Lowpass|Add3~38\);

-- Location: LABCELL_X33_Y65_N27
\TheRxFsk|Lowpass|Add3~33\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add3~33_sumout\ = SUM(( GND ) + ( \TheRxFsk|Lowpass|Mult0~32\ ) + ( \TheRxFsk|Lowpass|Add3~38\ ))
-- \TheRxFsk|Lowpass|Add3~34\ = CARRY(( GND ) + ( \TheRxFsk|Lowpass|Mult0~32\ ) + ( \TheRxFsk|Lowpass|Add3~38\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Lowpass|ALT_INV_Mult0~32\,
	cin => \TheRxFsk|Lowpass|Add3~38\,
	sumout => \TheRxFsk|Lowpass|Add3~33_sumout\,
	cout => \TheRxFsk|Lowpass|Add3~34\);

-- Location: LABCELL_X33_Y65_N30
\TheRxFsk|Lowpass|Add3~29\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add3~29_sumout\ = SUM(( GND ) + ( \TheRxFsk|Lowpass|Mult0~33\ ) + ( \TheRxFsk|Lowpass|Add3~34\ ))
-- \TheRxFsk|Lowpass|Add3~30\ = CARRY(( GND ) + ( \TheRxFsk|Lowpass|Mult0~33\ ) + ( \TheRxFsk|Lowpass|Add3~34\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Lowpass|ALT_INV_Mult0~33\,
	cin => \TheRxFsk|Lowpass|Add3~34\,
	sumout => \TheRxFsk|Lowpass|Add3~29_sumout\,
	cout => \TheRxFsk|Lowpass|Add3~30\);

-- Location: LABCELL_X33_Y65_N33
\TheRxFsk|Lowpass|Add3~25\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add3~25_sumout\ = SUM(( GND ) + ( \TheRxFsk|Lowpass|Mult0~34\ ) + ( \TheRxFsk|Lowpass|Add3~30\ ))
-- \TheRxFsk|Lowpass|Add3~26\ = CARRY(( GND ) + ( \TheRxFsk|Lowpass|Mult0~34\ ) + ( \TheRxFsk|Lowpass|Add3~30\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Lowpass|ALT_INV_Mult0~34\,
	cin => \TheRxFsk|Lowpass|Add3~30\,
	sumout => \TheRxFsk|Lowpass|Add3~25_sumout\,
	cout => \TheRxFsk|Lowpass|Add3~26\);

-- Location: LABCELL_X33_Y65_N36
\TheRxFsk|Lowpass|Add3~21\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add3~21_sumout\ = SUM(( \TheRxFsk|Lowpass|Mult0~35\ ) + ( GND ) + ( \TheRxFsk|Lowpass|Add3~26\ ))
-- \TheRxFsk|Lowpass|Add3~22\ = CARRY(( \TheRxFsk|Lowpass|Mult0~35\ ) + ( GND ) + ( \TheRxFsk|Lowpass|Add3~26\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datad => \TheRxFsk|Lowpass|ALT_INV_Mult0~35\,
	cin => \TheRxFsk|Lowpass|Add3~26\,
	sumout => \TheRxFsk|Lowpass|Add3~21_sumout\,
	cout => \TheRxFsk|Lowpass|Add3~22\);

-- Location: LABCELL_X33_Y65_N39
\TheRxFsk|Lowpass|Add3~17\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add3~17_sumout\ = SUM(( GND ) + ( \TheRxFsk|Lowpass|Mult0~36\ ) + ( \TheRxFsk|Lowpass|Add3~22\ ))
-- \TheRxFsk|Lowpass|Add3~18\ = CARRY(( GND ) + ( \TheRxFsk|Lowpass|Mult0~36\ ) + ( \TheRxFsk|Lowpass|Add3~22\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Lowpass|ALT_INV_Mult0~36\,
	cin => \TheRxFsk|Lowpass|Add3~22\,
	sumout => \TheRxFsk|Lowpass|Add3~17_sumout\,
	cout => \TheRxFsk|Lowpass|Add3~18\);

-- Location: LABCELL_X33_Y65_N42
\TheRxFsk|Lowpass|Add3~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add3~13_sumout\ = SUM(( GND ) + ( \TheRxFsk|Lowpass|Mult0~37\ ) + ( \TheRxFsk|Lowpass|Add3~18\ ))
-- \TheRxFsk|Lowpass|Add3~14\ = CARRY(( GND ) + ( \TheRxFsk|Lowpass|Mult0~37\ ) + ( \TheRxFsk|Lowpass|Add3~18\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Lowpass|ALT_INV_Mult0~37\,
	cin => \TheRxFsk|Lowpass|Add3~18\,
	sumout => \TheRxFsk|Lowpass|Add3~13_sumout\,
	cout => \TheRxFsk|Lowpass|Add3~14\);

-- Location: LABCELL_X33_Y65_N45
\TheRxFsk|Lowpass|Add3~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add3~9_sumout\ = SUM(( GND ) + ( \TheRxFsk|Lowpass|Mult0~38\ ) + ( \TheRxFsk|Lowpass|Add3~14\ ))
-- \TheRxFsk|Lowpass|Add3~10\ = CARRY(( GND ) + ( \TheRxFsk|Lowpass|Mult0~38\ ) + ( \TheRxFsk|Lowpass|Add3~14\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Lowpass|ALT_INV_Mult0~38\,
	cin => \TheRxFsk|Lowpass|Add3~14\,
	sumout => \TheRxFsk|Lowpass|Add3~9_sumout\,
	cout => \TheRxFsk|Lowpass|Add3~10\);

-- Location: LABCELL_X33_Y65_N48
\TheRxFsk|Lowpass|Add3~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add3~5_sumout\ = SUM(( GND ) + ( \TheRxFsk|Lowpass|Mult0~39\ ) + ( \TheRxFsk|Lowpass|Add3~10\ ))
-- \TheRxFsk|Lowpass|Add3~6\ = CARRY(( GND ) + ( \TheRxFsk|Lowpass|Mult0~39\ ) + ( \TheRxFsk|Lowpass|Add3~10\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Lowpass|ALT_INV_Mult0~39\,
	cin => \TheRxFsk|Lowpass|Add3~10\,
	sumout => \TheRxFsk|Lowpass|Add3~5_sumout\,
	cout => \TheRxFsk|Lowpass|Add3~6\);

-- Location: LABCELL_X33_Y65_N51
\TheRxFsk|Lowpass|Add3~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add3~1_sumout\ = SUM(( VCC ) + ( \TheRxFsk|Lowpass|Mult0~39\ ) + ( \TheRxFsk|Lowpass|Add3~6\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000101010101010101000000000000000001111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_Mult0~39\,
	cin => \TheRxFsk|Lowpass|Add3~6\,
	sumout => \TheRxFsk|Lowpass|Add3~1_sumout\);

-- Location: MLABCELL_X34_Y64_N36
\TheRxFsk|Lowpass|MultResultDelayed[0]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|MultResultDelayed[0]~0_combout\ = ( !\TheRxFsk|Lowpass|Add3~1_sumout\ )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111111111111111111111111111100000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \TheRxFsk|Lowpass|ALT_INV_Add3~1_sumout\,
	combout => \TheRxFsk|Lowpass|MultResultDelayed[0]~0_combout\);

-- Location: FF_X34_Y64_N37
\TheRxFsk|Lowpass|MultResultDelayed[0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|MultResultDelayed[0]~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|MultResultDelayed\(0));

-- Location: FF_X33_Y65_N46
\TheRxFsk|Lowpass|MultResultDelayed[-15]_NEW_REG4\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|Add3~9_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM5\);

-- Location: FF_X33_Y65_N43
\TheRxFsk|Lowpass|MultResultDelayed[-1]_NEW_REG18\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|Add3~13_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|MultResultDelayed[-1]_OTERM19\);

-- Location: FF_X33_Y65_N53
\TheRxFsk|Lowpass|MultResultDelayed[-15]_NEW_REG0\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|Add3~1_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM1\);

-- Location: FF_X33_Y65_N49
\TheRxFsk|Lowpass|MultResultDelayed[-15]_NEW_REG2\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|Add3~5_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM3\);

-- Location: MLABCELL_X34_Y65_N0
\TheRxFsk|Lowpass|MultResult[-1]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|MultResult[-1]~0_combout\ = ( \TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM3\ & ( ((\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM5\ & \TheRxFsk|Lowpass|MultResultDelayed[-1]_OTERM19\)) # 
-- (\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM1\) ) ) # ( !\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM3\ & ( (\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM1\ & ((\TheRxFsk|Lowpass|MultResultDelayed[-1]_OTERM19\) # 
-- (\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM5\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000011100000111000111110001111100000111000001110001111100011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM5\,
	datab => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-1]_OTERM19\,
	datac => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM1\,
	datae => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM3\,
	combout => \TheRxFsk|Lowpass|MultResult[-1]~0_combout\);

-- Location: LABCELL_X31_Y62_N45
\TheRxFsk|Lowpass|Add4~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add4~5_sumout\ = SUM(( \TheRxFsk|Lowpass|Sum\(0) ) + ( \TheRxFsk|Lowpass|MultResultDelayed\(0) ) + ( \TheRxFsk|Lowpass|Add4~10\ ))
-- \TheRxFsk|Lowpass|Add4~6\ = CARRY(( \TheRxFsk|Lowpass|Sum\(0) ) + ( \TheRxFsk|Lowpass|MultResultDelayed\(0) ) + ( \TheRxFsk|Lowpass|Add4~10\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111110000000000000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Lowpass|ALT_INV_Sum\(0),
	dataf => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed\(0),
	cin => \TheRxFsk|Lowpass|Add4~10\,
	sumout => \TheRxFsk|Lowpass|Add4~5_sumout\,
	cout => \TheRxFsk|Lowpass|Add4~6\);

-- Location: FF_X33_Y65_N40
\TheRxFsk|Lowpass|MultResultDelayed[-2]_NEW_REG22\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|Add3~17_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|MultResultDelayed[-2]_OTERM23\);

-- Location: MLABCELL_X34_Y65_N54
\TheRxFsk|Lowpass|MultResult[-2]~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|MultResult[-2]~1_combout\ = ( \TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM3\ & ( \TheRxFsk|Lowpass|MultResultDelayed[-2]_OTERM23\ & ( (\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM1\) # 
-- (\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM5\) ) ) ) # ( !\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM3\ & ( \TheRxFsk|Lowpass|MultResultDelayed[-2]_OTERM23\ & ( \TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM1\ ) ) ) # ( 
-- \TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM3\ & ( !\TheRxFsk|Lowpass|MultResultDelayed[-2]_OTERM23\ & ( \TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM1\ ) ) ) # ( !\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM3\ & ( 
-- !\TheRxFsk|Lowpass|MultResultDelayed[-2]_OTERM23\ & ( (\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM5\ & \TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM1\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100000101000011110000111100001111000011110101111101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM5\,
	datac => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM1\,
	datae => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM3\,
	dataf => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-2]_OTERM23\,
	combout => \TheRxFsk|Lowpass|MultResult[-2]~1_combout\);

-- Location: FF_X33_Y65_N37
\TheRxFsk|Lowpass|MultResultDelayed[-3]_NEW_REG26\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|Add3~21_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|MultResultDelayed[-3]_OTERM27\);

-- Location: MLABCELL_X34_Y65_N51
\TheRxFsk|Lowpass|MultResult[-3]~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|MultResult[-3]~2_combout\ = ( \TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM3\ & ( \TheRxFsk|Lowpass|MultResultDelayed[-3]_OTERM27\ & ( (\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM5\) # 
-- (\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM1\) ) ) ) # ( !\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM3\ & ( \TheRxFsk|Lowpass|MultResultDelayed[-3]_OTERM27\ & ( \TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM1\ ) ) ) # ( 
-- \TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM3\ & ( !\TheRxFsk|Lowpass|MultResultDelayed[-3]_OTERM27\ & ( \TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM1\ ) ) ) # ( !\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM3\ & ( 
-- !\TheRxFsk|Lowpass|MultResultDelayed[-3]_OTERM27\ & ( (\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM1\ & \TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM5\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001010101010101010101010101010101010101010101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM1\,
	datad => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM5\,
	datae => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM3\,
	dataf => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-3]_OTERM27\,
	combout => \TheRxFsk|Lowpass|MultResult[-3]~2_combout\);

-- Location: FF_X33_Y65_N34
\TheRxFsk|Lowpass|MultResultDelayed[-4]_NEW_REG30\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|Add3~25_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|MultResultDelayed[-4]_OTERM31\);

-- Location: MLABCELL_X34_Y65_N6
\TheRxFsk|Lowpass|MultResult[-4]~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|MultResult[-4]~3_combout\ = ( \TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM3\ & ( ((\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM5\ & \TheRxFsk|Lowpass|MultResultDelayed[-4]_OTERM31\)) # 
-- (\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM1\) ) ) # ( !\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM3\ & ( (\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM1\ & ((\TheRxFsk|Lowpass|MultResultDelayed[-4]_OTERM31\) # 
-- (\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM5\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000011100000111000111110001111100000111000001110001111100011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM5\,
	datab => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-4]_OTERM31\,
	datac => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM1\,
	datae => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM3\,
	combout => \TheRxFsk|Lowpass|MultResult[-4]~3_combout\);

-- Location: FF_X33_Y65_N31
\TheRxFsk|Lowpass|MultResultDelayed[-5]_NEW_REG34\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|Add3~29_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|MultResultDelayed[-5]_OTERM35\);

-- Location: MLABCELL_X34_Y65_N39
\TheRxFsk|Lowpass|MultResult[-5]~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|MultResult[-5]~4_combout\ = ( \TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM3\ & ( \TheRxFsk|Lowpass|MultResultDelayed[-5]_OTERM35\ & ( (\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM5\) # 
-- (\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM1\) ) ) ) # ( !\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM3\ & ( \TheRxFsk|Lowpass|MultResultDelayed[-5]_OTERM35\ & ( \TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM1\ ) ) ) # ( 
-- \TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM3\ & ( !\TheRxFsk|Lowpass|MultResultDelayed[-5]_OTERM35\ & ( \TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM1\ ) ) ) # ( !\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM3\ & ( 
-- !\TheRxFsk|Lowpass|MultResultDelayed[-5]_OTERM35\ & ( (\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM1\ & \TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM5\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000001010101010101010101010101010101010101010101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM1\,
	datad => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM5\,
	datae => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM3\,
	dataf => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-5]_OTERM35\,
	combout => \TheRxFsk|Lowpass|MultResult[-5]~4_combout\);

-- Location: FF_X33_Y65_N28
\TheRxFsk|Lowpass|MultResultDelayed[-6]_NEW_REG38\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|Add3~33_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|MultResultDelayed[-6]_OTERM39\);

-- Location: MLABCELL_X34_Y65_N42
\TheRxFsk|Lowpass|MultResult[-6]~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|MultResult[-6]~5_combout\ = ( \TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM1\ & ( ((\TheRxFsk|Lowpass|MultResultDelayed[-6]_OTERM39\) # (\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM3\)) # 
-- (\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM5\) ) ) # ( !\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM1\ & ( (\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM5\ & (\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM3\ & 
-- \TheRxFsk|Lowpass|MultResultDelayed[-6]_OTERM39\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000100000001000000010000000101111111011111110111111101111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM5\,
	datab => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM3\,
	datac => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-6]_OTERM39\,
	dataf => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM1\,
	combout => \TheRxFsk|Lowpass|MultResult[-6]~5_combout\);

-- Location: FF_X33_Y65_N25
\TheRxFsk|Lowpass|MultResultDelayed[-7]_NEW_REG40\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|Add3~37_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|MultResultDelayed[-7]_OTERM41\);

-- Location: MLABCELL_X34_Y65_N45
\TheRxFsk|Lowpass|MultResult[-7]~6\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|MultResult[-7]~6_combout\ = ( \TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM1\ & ( ((\TheRxFsk|Lowpass|MultResultDelayed[-7]_OTERM41\) # (\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM3\)) # 
-- (\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM5\) ) ) # ( !\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM1\ & ( (\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM5\ & (\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM3\ & 
-- \TheRxFsk|Lowpass|MultResultDelayed[-7]_OTERM41\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000100000001000000010000000101111111011111110111111101111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM5\,
	datab => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM3\,
	datac => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-7]_OTERM41\,
	dataf => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM1\,
	combout => \TheRxFsk|Lowpass|MultResult[-7]~6_combout\);

-- Location: FF_X33_Y65_N22
\TheRxFsk|Lowpass|MultResultDelayed[-8]_NEW_REG44\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|Add3~41_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|MultResultDelayed[-8]_OTERM45\);

-- Location: MLABCELL_X34_Y65_N12
\TheRxFsk|Lowpass|MultResult[-8]~7\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|MultResult[-8]~7_combout\ = ( \TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM1\ & ( ((\TheRxFsk|Lowpass|MultResultDelayed[-8]_OTERM45\) # (\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM3\)) # 
-- (\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM5\) ) ) # ( !\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM1\ & ( (\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM5\ & (\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM3\ & 
-- \TheRxFsk|Lowpass|MultResultDelayed[-8]_OTERM45\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000100000001000000010000000101111111011111110111111101111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM5\,
	datab => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM3\,
	datac => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-8]_OTERM45\,
	dataf => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM1\,
	combout => \TheRxFsk|Lowpass|MultResult[-8]~7_combout\);

-- Location: FF_X33_Y65_N19
\TheRxFsk|Lowpass|MultResultDelayed[-9]_NEW_REG50\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|Add3~45_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|MultResultDelayed[-9]_OTERM51\);

-- Location: MLABCELL_X34_Y65_N15
\TheRxFsk|Lowpass|MultResult[-9]~8\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|MultResult[-9]~8_combout\ = ( \TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM1\ & ( ((\TheRxFsk|Lowpass|MultResultDelayed[-9]_OTERM51\) # (\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM3\)) # 
-- (\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM5\) ) ) # ( !\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM1\ & ( (\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM5\ & (\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM3\ & 
-- \TheRxFsk|Lowpass|MultResultDelayed[-9]_OTERM51\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000100000001000000010000000101111111011111110111111101111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM5\,
	datab => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM3\,
	datac => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-9]_OTERM51\,
	dataf => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM1\,
	combout => \TheRxFsk|Lowpass|MultResult[-9]~8_combout\);

-- Location: FF_X33_Y65_N16
\TheRxFsk|Lowpass|MultResultDelayed[-10]_NEW_REG48\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|Add3~49_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|MultResultDelayed[-10]_OTERM49\);

-- Location: MLABCELL_X34_Y65_N21
\TheRxFsk|Lowpass|MultResult[-10]~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|MultResult[-10]~9_combout\ = ( \TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM3\ & ( \TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM5\ & ( (\TheRxFsk|Lowpass|MultResultDelayed[-10]_OTERM49\) # 
-- (\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM1\) ) ) ) # ( !\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM3\ & ( \TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM5\ & ( \TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM1\ ) ) ) # ( 
-- \TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM3\ & ( !\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM5\ & ( \TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM1\ ) ) ) # ( !\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM3\ & ( 
-- !\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM5\ & ( (\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM1\ & \TheRxFsk|Lowpass|MultResultDelayed[-10]_OTERM49\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010100000101010101010101010101010101010101010101111101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM1\,
	datac => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-10]_OTERM49\,
	datae => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM3\,
	dataf => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM5\,
	combout => \TheRxFsk|Lowpass|MultResult[-10]~9_combout\);

-- Location: FF_X33_Y65_N13
\TheRxFsk|Lowpass|MultResultDelayed[-11]_NEW_REG56\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|Add3~53_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|MultResultDelayed[-11]_OTERM57\);

-- Location: MLABCELL_X34_Y65_N24
\TheRxFsk|Lowpass|MultResult[-11]~10\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|MultResult[-11]~10_combout\ = ( \TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM1\ & ( ((\TheRxFsk|Lowpass|MultResultDelayed[-11]_OTERM57\) # (\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM3\)) # 
-- (\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM5\) ) ) # ( !\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM1\ & ( (\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM5\ & (\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM3\ & 
-- \TheRxFsk|Lowpass|MultResultDelayed[-11]_OTERM57\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000100000001000000010000000101111111011111110111111101111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM5\,
	datab => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM3\,
	datac => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-11]_OTERM57\,
	dataf => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM1\,
	combout => \TheRxFsk|Lowpass|MultResult[-11]~10_combout\);

-- Location: FF_X33_Y65_N10
\TheRxFsk|Lowpass|MultResultDelayed[-12]_NEW_REG60\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|Add3~57_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|MultResultDelayed[-12]_OTERM61\);

-- Location: MLABCELL_X34_Y65_N27
\TheRxFsk|Lowpass|MultResult[-12]~11\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|MultResult[-12]~11_combout\ = ( \TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM1\ & ( ((\TheRxFsk|Lowpass|MultResultDelayed[-12]_OTERM61\) # (\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM3\)) # 
-- (\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM5\) ) ) # ( !\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM1\ & ( (\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM5\ & (\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM3\ & 
-- \TheRxFsk|Lowpass|MultResultDelayed[-12]_OTERM61\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000100000001000000010000000101111111011111110111111101111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM5\,
	datab => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM3\,
	datac => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-12]_OTERM61\,
	dataf => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM1\,
	combout => \TheRxFsk|Lowpass|MultResult[-12]~11_combout\);

-- Location: FF_X33_Y65_N7
\TheRxFsk|Lowpass|MultResultDelayed[-13]_NEW_REG88\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|Add3~61_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|MultResultDelayed[-13]_OTERM89\);

-- Location: MLABCELL_X34_Y65_N30
\TheRxFsk|Lowpass|MultResult[-13]~12\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|MultResult[-13]~12_combout\ = ( \TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM1\ & ( ((\TheRxFsk|Lowpass|MultResultDelayed[-13]_OTERM89\) # (\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM3\)) # 
-- (\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM5\) ) ) # ( !\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM1\ & ( (\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM5\ & (\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM3\ & 
-- \TheRxFsk|Lowpass|MultResultDelayed[-13]_OTERM89\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000100000001000000010000000101111111011111110111111101111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM5\,
	datab => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM3\,
	datac => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-13]_OTERM89\,
	dataf => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM1\,
	combout => \TheRxFsk|Lowpass|MultResult[-13]~12_combout\);

-- Location: FF_X33_Y65_N4
\TheRxFsk|Lowpass|MultResultDelayed[-14]_NEW_REG92\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|Add3~65_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|MultResultDelayed[-14]_OTERM93\);

-- Location: MLABCELL_X34_Y65_N33
\TheRxFsk|Lowpass|MultResult[-14]~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|MultResult[-14]~13_combout\ = ( \TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM1\ & ( ((\TheRxFsk|Lowpass|MultResultDelayed[-14]_OTERM93\) # (\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM3\)) # 
-- (\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM5\) ) ) # ( !\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM1\ & ( (\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM5\ & (\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM3\ & 
-- \TheRxFsk|Lowpass|MultResultDelayed[-14]_OTERM93\)) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000100000001000000010000000101111111011111110111111101111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM5\,
	datab => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM3\,
	datac => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-14]_OTERM93\,
	dataf => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM1\,
	combout => \TheRxFsk|Lowpass|MultResult[-14]~13_combout\);

-- Location: FF_X33_Y65_N1
\TheRxFsk|Lowpass|MultResultDelayed[-15]_NEW_REG6\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|Add3~69_sumout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM7\);

-- Location: MLABCELL_X34_Y62_N39
\TheRxFsk|Lowpass|MultResult[-15]~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|MultResult[-15]~14_combout\ = ( \TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM7\ & ( ((\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM3\ & \TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM5\)) # 
-- (\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM1\) ) ) # ( !\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM7\ & ( (\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM1\ & ((\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM5\) # 
-- (\TheRxFsk|Lowpass|MultResultDelayed[-15]_OTERM3\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100001111000000110000111100001111001111110000111100111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM3\,
	datac => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM1\,
	datad => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM5\,
	dataf => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed[-15]_OTERM7\,
	combout => \TheRxFsk|Lowpass|MultResult[-15]~14_combout\);

-- Location: LABCELL_X30_Y62_N54
\TheRxFsk|Lowpass|NextSum[-15]~14\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|NextSum[-15]~14_combout\ = ( \TheRxFsk|Lowpass|Sum[-15]~q\ & ( \TheRxFsk|Lowpass|MultResult[-15]~14_combout\ & ( (\TheRxFsk|Lowpass|Add4~1_sumout\ & \TheRxFsk|Lowpass|Add4~5_sumout\) ) ) ) # ( !\TheRxFsk|Lowpass|Sum[-15]~q\ & ( 
-- \TheRxFsk|Lowpass|MultResult[-15]~14_combout\ & ( (\TheRxFsk|Lowpass|Add4~5_sumout\) # (\TheRxFsk|Lowpass|Add4~1_sumout\) ) ) ) # ( \TheRxFsk|Lowpass|Sum[-15]~q\ & ( !\TheRxFsk|Lowpass|MultResult[-15]~14_combout\ & ( (\TheRxFsk|Lowpass|Add4~5_sumout\) # 
-- (\TheRxFsk|Lowpass|Add4~1_sumout\) ) ) ) # ( !\TheRxFsk|Lowpass|Sum[-15]~q\ & ( !\TheRxFsk|Lowpass|MultResult[-15]~14_combout\ & ( (\TheRxFsk|Lowpass|Add4~1_sumout\ & \TheRxFsk|Lowpass|Add4~5_sumout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000001100000011001111110011111100111111001111110000001100000011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Lowpass|ALT_INV_Add4~1_sumout\,
	datac => \TheRxFsk|Lowpass|ALT_INV_Add4~5_sumout\,
	datae => \TheRxFsk|Lowpass|ALT_INV_Sum[-15]~q\,
	dataf => \TheRxFsk|Lowpass|ALT_INV_MultResult[-15]~14_combout\,
	combout => \TheRxFsk|Lowpass|NextSum[-15]~14_combout\);

-- Location: FF_X31_Y62_N52
\TheRxFsk|Lowpass|R.SumState.SumValid\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	asdata => \TheRxFsk|Lowpass|R.SumState.SumWait2~DUPLICATE_q\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|R.SumState.SumValid~q\);

-- Location: LABCELL_X29_Y62_N48
\TheRxFsk|Lowpass|Selector0~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Selector0~0_combout\ = ( \TheRxFsk|Lowpass|R.SumState.Idle~q\ & ( !\TheRxFsk|Lowpass|R.SumState.SumValid~q\ ) ) # ( !\TheRxFsk|Lowpass|R.SumState.Idle~q\ & ( (\TheRxFsk|Bandpasses:11:Bandpass0|R.ValWet~q\ & 
-- !\TheRxFsk|Lowpass|R.SumState.SumValid~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100000000111111110000000000001111000000001111111100000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Bandpasses:11:Bandpass0|ALT_INV_R.ValWet~q\,
	datad => \TheRxFsk|Lowpass|ALT_INV_R.SumState.SumValid~q\,
	datae => \TheRxFsk|Lowpass|ALT_INV_R.SumState.Idle~q\,
	combout => \TheRxFsk|Lowpass|Selector0~0_combout\);

-- Location: FF_X29_Y62_N50
\TheRxFsk|Lowpass|R.SumState.Idle\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|Selector0~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|R.SumState.Idle~q\);

-- Location: LABCELL_X29_Y62_N45
\TheRxFsk|Lowpass|Selector1~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Selector1~0_combout\ = ( \TheRxFsk|Bandpasses:11:Bandpass0|R.ValWet~q\ & ( !\TheRxFsk|Lowpass|R.SumState.Idle~q\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111111111111100000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datae => \TheRxFsk|Bandpasses:11:Bandpass0|ALT_INV_R.ValWet~q\,
	dataf => \TheRxFsk|Lowpass|ALT_INV_R.SumState.Idle~q\,
	combout => \TheRxFsk|Lowpass|Selector1~0_combout\);

-- Location: FF_X29_Y62_N46
\TheRxFsk|Lowpass|R.SumState.SumEnable\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|Selector1~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|R.SumState.SumEnable~q\);

-- Location: LABCELL_X29_Y62_N24
\TheRxFsk|Lowpass|Selector2~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Selector2~0_combout\ = ( \TheRxFsk|Lowpass|R.SumState.SumEnable~q\ ) # ( !\TheRxFsk|Lowpass|R.SumState.SumEnable~q\ & ( (\TheRxFsk|Lowpass|R.SumState.SumSelect~q\ & ((!\TheRxFsk|Lowpass|CoefMemory~0_combout\) # 
-- (!\TheRxFsk|Lowpass|Equal1~0_combout\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011101110000000001110111011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_CoefMemory~0_combout\,
	datab => \TheRxFsk|Lowpass|ALT_INV_Equal1~0_combout\,
	datad => \TheRxFsk|Lowpass|ALT_INV_R.SumState.SumSelect~q\,
	dataf => \TheRxFsk|Lowpass|ALT_INV_R.SumState.SumEnable~q\,
	combout => \TheRxFsk|Lowpass|Selector2~0_combout\);

-- Location: FF_X29_Y62_N25
\TheRxFsk|Lowpass|R.SumState.SumSelect\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|Selector2~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|R.SumState.SumSelect~q\);

-- Location: LABCELL_X29_Y62_N27
\TheRxFsk|Lowpass|Selector3~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Selector3~0_combout\ = ( \TheRxFsk|Lowpass|R.SumState.SumSelect~q\ & ( (\TheRxFsk|Lowpass|CoefMemory~0_combout\ & \TheRxFsk|Lowpass|Equal1~0_combout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000010001000100010001000100010001",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_CoefMemory~0_combout\,
	datab => \TheRxFsk|Lowpass|ALT_INV_Equal1~0_combout\,
	dataf => \TheRxFsk|Lowpass|ALT_INV_R.SumState.SumSelect~q\,
	combout => \TheRxFsk|Lowpass|Selector3~0_combout\);

-- Location: FF_X29_Y62_N29
\TheRxFsk|Lowpass|R.SumState.SumWait1\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|Selector3~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|R.SumState.SumWait1~q\);

-- Location: FF_X29_Y62_N16
\TheRxFsk|Lowpass|R.SumState.SumWait2~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	asdata => \TheRxFsk|Lowpass|R.SumState.SumWait1~q\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|R.SumState.SumWait2~DUPLICATE_q\);

-- Location: LABCELL_X31_Y62_N54
\TheRxFsk|Lowpass|Selector6~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Selector6~0_combout\ = ( \TheRxFsk|Lowpass|R.SelSumUp~q\ & ( \TheRxFsk|Lowpass|R.SumState.SumEnable~q\ ) ) # ( !\TheRxFsk|Lowpass|R.SelSumUp~q\ & ( \TheRxFsk|Lowpass|R.SumState.SumEnable~q\ ) ) # ( \TheRxFsk|Lowpass|R.SelSumUp~q\ & ( 
-- !\TheRxFsk|Lowpass|R.SumState.SumEnable~q\ & ( !\TheRxFsk|Lowpass|R.SumState.SumWait2~DUPLICATE_q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000101010101010101011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_R.SumState.SumWait2~DUPLICATE_q\,
	datae => \TheRxFsk|Lowpass|ALT_INV_R.SelSumUp~q\,
	dataf => \TheRxFsk|Lowpass|ALT_INV_R.SumState.SumEnable~q\,
	combout => \TheRxFsk|Lowpass|Selector6~0_combout\);

-- Location: FF_X31_Y62_N56
\TheRxFsk|Lowpass|R.SelSumUp\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|Selector6~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|R.SelSumUp~q\);

-- Location: FF_X29_Y62_N17
\TheRxFsk|Lowpass|R.SumState.SumWait2\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	asdata => \TheRxFsk|Lowpass|R.SumState.SumWait1~q\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => VCC,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|R.SumState.SumWait2~q\);

-- Location: LABCELL_X29_Y62_N21
\TheRxFsk|Lowpass|Selector7~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Selector7~0_combout\ = ( \TheRxFsk|Lowpass|R.EnableSumUp~q\ & ( \TheRxFsk|Lowpass|R.SumState.Idle~q\ & ( !\TheRxFsk|Lowpass|R.SumState.SumWait2~q\ ) ) ) # ( \TheRxFsk|Lowpass|R.EnableSumUp~q\ & ( !\TheRxFsk|Lowpass|R.SumState.Idle~q\ ) ) 
-- # ( !\TheRxFsk|Lowpass|R.EnableSumUp~q\ & ( !\TheRxFsk|Lowpass|R.SumState.Idle~q\ & ( \TheRxFsk|Bandpasses:11:Bandpass0|R.ValWet~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010101010101111111111111111100000000000000001100110011001100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Bandpasses:11:Bandpass0|ALT_INV_R.ValWet~q\,
	datab => \TheRxFsk|Lowpass|ALT_INV_R.SumState.SumWait2~q\,
	datae => \TheRxFsk|Lowpass|ALT_INV_R.EnableSumUp~q\,
	dataf => \TheRxFsk|Lowpass|ALT_INV_R.SumState.Idle~q\,
	combout => \TheRxFsk|Lowpass|Selector7~0_combout\);

-- Location: FF_X29_Y62_N22
\TheRxFsk|Lowpass|R.EnableSumUp\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|Selector7~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|R.EnableSumUp~q\);

-- Location: FF_X30_Y62_N55
\TheRxFsk|Lowpass|Sum[-15]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|NextSum[-15]~14_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Lowpass|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Lowpass|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|Sum[-15]~q\);

-- Location: LABCELL_X31_Y62_N0
\TheRxFsk|Lowpass|Add4~65\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add4~66\ = CARRY(( \TheRxFsk|Lowpass|MultResult[-15]~14_combout\ ) + ( \TheRxFsk|Lowpass|Sum[-15]~q\ ) + ( !VCC ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111110000000000000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Lowpass|ALT_INV_MultResult[-15]~14_combout\,
	dataf => \TheRxFsk|Lowpass|ALT_INV_Sum[-15]~q\,
	cin => GND,
	cout => \TheRxFsk|Lowpass|Add4~66\);

-- Location: LABCELL_X31_Y62_N3
\TheRxFsk|Lowpass|Add4~61\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add4~61_sumout\ = SUM(( \TheRxFsk|Lowpass|Sum[-14]~q\ ) + ( \TheRxFsk|Lowpass|MultResult[-14]~13_combout\ ) + ( \TheRxFsk|Lowpass|Add4~66\ ))
-- \TheRxFsk|Lowpass|Add4~62\ = CARRY(( \TheRxFsk|Lowpass|Sum[-14]~q\ ) + ( \TheRxFsk|Lowpass|MultResult[-14]~13_combout\ ) + ( \TheRxFsk|Lowpass|Add4~66\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000101010101010101000000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_MultResult[-14]~13_combout\,
	datac => \TheRxFsk|Lowpass|ALT_INV_Sum[-14]~q\,
	cin => \TheRxFsk|Lowpass|Add4~66\,
	sumout => \TheRxFsk|Lowpass|Add4~61_sumout\,
	cout => \TheRxFsk|Lowpass|Add4~62\);

-- Location: LABCELL_X30_Y62_N15
\TheRxFsk|Lowpass|NextSum[-14]~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|NextSum[-14]~13_combout\ = (!\TheRxFsk|Lowpass|Add4~5_sumout\ & (\TheRxFsk|Lowpass|Add4~1_sumout\ & \TheRxFsk|Lowpass|Add4~61_sumout\)) # (\TheRxFsk|Lowpass|Add4~5_sumout\ & ((\TheRxFsk|Lowpass|Add4~61_sumout\) # 
-- (\TheRxFsk|Lowpass|Add4~1_sumout\)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000101110111000100010111011100010001011101110001000101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_Add4~5_sumout\,
	datab => \TheRxFsk|Lowpass|ALT_INV_Add4~1_sumout\,
	datad => \TheRxFsk|Lowpass|ALT_INV_Add4~61_sumout\,
	combout => \TheRxFsk|Lowpass|NextSum[-14]~13_combout\);

-- Location: FF_X30_Y62_N16
\TheRxFsk|Lowpass|Sum[-14]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|NextSum[-14]~13_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Lowpass|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Lowpass|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|Sum[-14]~q\);

-- Location: LABCELL_X31_Y62_N6
\TheRxFsk|Lowpass|Add4~57\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add4~57_sumout\ = SUM(( \TheRxFsk|Lowpass|Sum[-13]~q\ ) + ( \TheRxFsk|Lowpass|MultResult[-13]~12_combout\ ) + ( \TheRxFsk|Lowpass|Add4~62\ ))
-- \TheRxFsk|Lowpass|Add4~58\ = CARRY(( \TheRxFsk|Lowpass|Sum[-13]~q\ ) + ( \TheRxFsk|Lowpass|MultResult[-13]~12_combout\ ) + ( \TheRxFsk|Lowpass|Add4~62\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000101010101010101000000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_MultResult[-13]~12_combout\,
	datac => \TheRxFsk|Lowpass|ALT_INV_Sum[-13]~q\,
	cin => \TheRxFsk|Lowpass|Add4~62\,
	sumout => \TheRxFsk|Lowpass|Add4~57_sumout\,
	cout => \TheRxFsk|Lowpass|Add4~58\);

-- Location: LABCELL_X30_Y62_N12
\TheRxFsk|Lowpass|NextSum[-13]~12\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|NextSum[-13]~12_combout\ = (!\TheRxFsk|Lowpass|Add4~5_sumout\ & (\TheRxFsk|Lowpass|Add4~1_sumout\ & \TheRxFsk|Lowpass|Add4~57_sumout\)) # (\TheRxFsk|Lowpass|Add4~5_sumout\ & ((\TheRxFsk|Lowpass|Add4~57_sumout\) # 
-- (\TheRxFsk|Lowpass|Add4~1_sumout\)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001011100010111000101110001011100010111000101110001011100010111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_Add4~5_sumout\,
	datab => \TheRxFsk|Lowpass|ALT_INV_Add4~1_sumout\,
	datac => \TheRxFsk|Lowpass|ALT_INV_Add4~57_sumout\,
	combout => \TheRxFsk|Lowpass|NextSum[-13]~12_combout\);

-- Location: FF_X30_Y62_N13
\TheRxFsk|Lowpass|Sum[-13]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|NextSum[-13]~12_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Lowpass|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Lowpass|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|Sum[-13]~q\);

-- Location: LABCELL_X31_Y62_N9
\TheRxFsk|Lowpass|Add4~53\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add4~53_sumout\ = SUM(( \TheRxFsk|Lowpass|MultResult[-12]~11_combout\ ) + ( \TheRxFsk|Lowpass|Sum[-12]~q\ ) + ( \TheRxFsk|Lowpass|Add4~58\ ))
-- \TheRxFsk|Lowpass|Add4~54\ = CARRY(( \TheRxFsk|Lowpass|MultResult[-12]~11_combout\ ) + ( \TheRxFsk|Lowpass|Sum[-12]~q\ ) + ( \TheRxFsk|Lowpass|Add4~58\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111110000000000000000000000000011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Lowpass|ALT_INV_MultResult[-12]~11_combout\,
	dataf => \TheRxFsk|Lowpass|ALT_INV_Sum[-12]~q\,
	cin => \TheRxFsk|Lowpass|Add4~58\,
	sumout => \TheRxFsk|Lowpass|Add4~53_sumout\,
	cout => \TheRxFsk|Lowpass|Add4~54\);

-- Location: LABCELL_X30_Y62_N45
\TheRxFsk|Lowpass|NextSum[-12]~11\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|NextSum[-12]~11_combout\ = (!\TheRxFsk|Lowpass|Add4~5_sumout\ & (\TheRxFsk|Lowpass|Add4~1_sumout\ & \TheRxFsk|Lowpass|Add4~53_sumout\)) # (\TheRxFsk|Lowpass|Add4~5_sumout\ & ((\TheRxFsk|Lowpass|Add4~53_sumout\) # 
-- (\TheRxFsk|Lowpass|Add4~1_sumout\)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000101110111000100010111011100010001011101110001000101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_Add4~5_sumout\,
	datab => \TheRxFsk|Lowpass|ALT_INV_Add4~1_sumout\,
	datad => \TheRxFsk|Lowpass|ALT_INV_Add4~53_sumout\,
	combout => \TheRxFsk|Lowpass|NextSum[-12]~11_combout\);

-- Location: FF_X30_Y62_N46
\TheRxFsk|Lowpass|Sum[-12]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|NextSum[-12]~11_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Lowpass|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Lowpass|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|Sum[-12]~q\);

-- Location: LABCELL_X31_Y62_N12
\TheRxFsk|Lowpass|Add4~49\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add4~49_sumout\ = SUM(( \TheRxFsk|Lowpass|MultResult[-11]~10_combout\ ) + ( \TheRxFsk|Lowpass|Sum[-11]~q\ ) + ( \TheRxFsk|Lowpass|Add4~54\ ))
-- \TheRxFsk|Lowpass|Add4~50\ = CARRY(( \TheRxFsk|Lowpass|MultResult[-11]~10_combout\ ) + ( \TheRxFsk|Lowpass|Sum[-11]~q\ ) + ( \TheRxFsk|Lowpass|Add4~54\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000110011001100110000000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Lowpass|ALT_INV_Sum[-11]~q\,
	datad => \TheRxFsk|Lowpass|ALT_INV_MultResult[-11]~10_combout\,
	cin => \TheRxFsk|Lowpass|Add4~54\,
	sumout => \TheRxFsk|Lowpass|Add4~49_sumout\,
	cout => \TheRxFsk|Lowpass|Add4~50\);

-- Location: LABCELL_X30_Y62_N42
\TheRxFsk|Lowpass|NextSum[-11]~10\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|NextSum[-11]~10_combout\ = ( \TheRxFsk|Lowpass|Add4~49_sumout\ & ( (\TheRxFsk|Lowpass|Add4~1_sumout\) # (\TheRxFsk|Lowpass|Add4~5_sumout\) ) ) # ( !\TheRxFsk|Lowpass|Add4~49_sumout\ & ( (\TheRxFsk|Lowpass|Add4~5_sumout\ & 
-- \TheRxFsk|Lowpass|Add4~1_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000100010001000100010001000101110111011101110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_Add4~5_sumout\,
	datab => \TheRxFsk|Lowpass|ALT_INV_Add4~1_sumout\,
	dataf => \TheRxFsk|Lowpass|ALT_INV_Add4~49_sumout\,
	combout => \TheRxFsk|Lowpass|NextSum[-11]~10_combout\);

-- Location: FF_X30_Y62_N43
\TheRxFsk|Lowpass|Sum[-11]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|NextSum[-11]~10_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Lowpass|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Lowpass|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|Sum[-11]~q\);

-- Location: LABCELL_X31_Y62_N15
\TheRxFsk|Lowpass|Add4~45\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add4~45_sumout\ = SUM(( \TheRxFsk|Lowpass|Sum[-10]~q\ ) + ( \TheRxFsk|Lowpass|MultResult[-10]~9_combout\ ) + ( \TheRxFsk|Lowpass|Add4~50\ ))
-- \TheRxFsk|Lowpass|Add4~46\ = CARRY(( \TheRxFsk|Lowpass|Sum[-10]~q\ ) + ( \TheRxFsk|Lowpass|MultResult[-10]~9_combout\ ) + ( \TheRxFsk|Lowpass|Add4~50\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000101010101010101000000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_MultResult[-10]~9_combout\,
	datac => \TheRxFsk|Lowpass|ALT_INV_Sum[-10]~q\,
	cin => \TheRxFsk|Lowpass|Add4~50\,
	sumout => \TheRxFsk|Lowpass|Add4~45_sumout\,
	cout => \TheRxFsk|Lowpass|Add4~46\);

-- Location: LABCELL_X30_Y62_N27
\TheRxFsk|Lowpass|NextSum[-10]~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|NextSum[-10]~9_combout\ = ( \TheRxFsk|Lowpass|Add4~45_sumout\ & ( \TheRxFsk|Lowpass|Add4~5_sumout\ ) ) # ( !\TheRxFsk|Lowpass|Add4~45_sumout\ & ( \TheRxFsk|Lowpass|Add4~5_sumout\ & ( \TheRxFsk|Lowpass|Add4~1_sumout\ ) ) ) # ( 
-- \TheRxFsk|Lowpass|Add4~45_sumout\ & ( !\TheRxFsk|Lowpass|Add4~5_sumout\ & ( \TheRxFsk|Lowpass|Add4~1_sumout\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000011110000111100001111000011111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Lowpass|ALT_INV_Add4~1_sumout\,
	datae => \TheRxFsk|Lowpass|ALT_INV_Add4~45_sumout\,
	dataf => \TheRxFsk|Lowpass|ALT_INV_Add4~5_sumout\,
	combout => \TheRxFsk|Lowpass|NextSum[-10]~9_combout\);

-- Location: FF_X30_Y62_N28
\TheRxFsk|Lowpass|Sum[-10]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|NextSum[-10]~9_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Lowpass|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Lowpass|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|Sum[-10]~q\);

-- Location: LABCELL_X31_Y62_N18
\TheRxFsk|Lowpass|Add4~41\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add4~41_sumout\ = SUM(( \TheRxFsk|Lowpass|Sum[-9]~q\ ) + ( \TheRxFsk|Lowpass|MultResult[-9]~8_combout\ ) + ( \TheRxFsk|Lowpass|Add4~46\ ))
-- \TheRxFsk|Lowpass|Add4~42\ = CARRY(( \TheRxFsk|Lowpass|Sum[-9]~q\ ) + ( \TheRxFsk|Lowpass|MultResult[-9]~8_combout\ ) + ( \TheRxFsk|Lowpass|Add4~46\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111100001111000000000000000000000011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Lowpass|ALT_INV_Sum[-9]~q\,
	datac => \TheRxFsk|Lowpass|ALT_INV_MultResult[-9]~8_combout\,
	cin => \TheRxFsk|Lowpass|Add4~46\,
	sumout => \TheRxFsk|Lowpass|Add4~41_sumout\,
	cout => \TheRxFsk|Lowpass|Add4~42\);

-- Location: LABCELL_X30_Y62_N9
\TheRxFsk|Lowpass|NextSum[-9]~8\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|NextSum[-9]~8_combout\ = (!\TheRxFsk|Lowpass|Add4~5_sumout\ & (\TheRxFsk|Lowpass|Add4~1_sumout\ & \TheRxFsk|Lowpass|Add4~41_sumout\)) # (\TheRxFsk|Lowpass|Add4~5_sumout\ & ((\TheRxFsk|Lowpass|Add4~41_sumout\) # 
-- (\TheRxFsk|Lowpass|Add4~1_sumout\)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001011100010111000101110001011100010111000101110001011100010111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_Add4~5_sumout\,
	datab => \TheRxFsk|Lowpass|ALT_INV_Add4~1_sumout\,
	datac => \TheRxFsk|Lowpass|ALT_INV_Add4~41_sumout\,
	combout => \TheRxFsk|Lowpass|NextSum[-9]~8_combout\);

-- Location: FF_X30_Y62_N10
\TheRxFsk|Lowpass|Sum[-9]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|NextSum[-9]~8_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Lowpass|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Lowpass|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|Sum[-9]~q\);

-- Location: LABCELL_X31_Y62_N21
\TheRxFsk|Lowpass|Add4~37\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add4~37_sumout\ = SUM(( \TheRxFsk|Lowpass|Sum[-8]~q\ ) + ( \TheRxFsk|Lowpass|MultResult[-8]~7_combout\ ) + ( \TheRxFsk|Lowpass|Add4~42\ ))
-- \TheRxFsk|Lowpass|Add4~38\ = CARRY(( \TheRxFsk|Lowpass|Sum[-8]~q\ ) + ( \TheRxFsk|Lowpass|MultResult[-8]~7_combout\ ) + ( \TheRxFsk|Lowpass|Add4~42\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000101010101010101000000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_MultResult[-8]~7_combout\,
	datad => \TheRxFsk|Lowpass|ALT_INV_Sum[-8]~q\,
	cin => \TheRxFsk|Lowpass|Add4~42\,
	sumout => \TheRxFsk|Lowpass|Add4~37_sumout\,
	cout => \TheRxFsk|Lowpass|Add4~38\);

-- Location: LABCELL_X30_Y62_N6
\TheRxFsk|Lowpass|NextSum[-8]~7\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|NextSum[-8]~7_combout\ = (!\TheRxFsk|Lowpass|Add4~5_sumout\ & (\TheRxFsk|Lowpass|Add4~1_sumout\ & \TheRxFsk|Lowpass|Add4~37_sumout\)) # (\TheRxFsk|Lowpass|Add4~5_sumout\ & ((\TheRxFsk|Lowpass|Add4~37_sumout\) # 
-- (\TheRxFsk|Lowpass|Add4~1_sumout\)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001011100010111000101110001011100010111000101110001011100010111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_Add4~5_sumout\,
	datab => \TheRxFsk|Lowpass|ALT_INV_Add4~1_sumout\,
	datac => \TheRxFsk|Lowpass|ALT_INV_Add4~37_sumout\,
	combout => \TheRxFsk|Lowpass|NextSum[-8]~7_combout\);

-- Location: FF_X30_Y62_N7
\TheRxFsk|Lowpass|Sum[-8]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|NextSum[-8]~7_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Lowpass|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Lowpass|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|Sum[-8]~q\);

-- Location: LABCELL_X31_Y62_N24
\TheRxFsk|Lowpass|Add4~33\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add4~33_sumout\ = SUM(( \TheRxFsk|Lowpass|Sum[-7]~q\ ) + ( \TheRxFsk|Lowpass|MultResult[-7]~6_combout\ ) + ( \TheRxFsk|Lowpass|Add4~38\ ))
-- \TheRxFsk|Lowpass|Add4~34\ = CARRY(( \TheRxFsk|Lowpass|Sum[-7]~q\ ) + ( \TheRxFsk|Lowpass|MultResult[-7]~6_combout\ ) + ( \TheRxFsk|Lowpass|Add4~38\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000110011001100110000000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Lowpass|ALT_INV_MultResult[-7]~6_combout\,
	datac => \TheRxFsk|Lowpass|ALT_INV_Sum[-7]~q\,
	cin => \TheRxFsk|Lowpass|Add4~38\,
	sumout => \TheRxFsk|Lowpass|Add4~33_sumout\,
	cout => \TheRxFsk|Lowpass|Add4~34\);

-- Location: LABCELL_X30_Y62_N51
\TheRxFsk|Lowpass|NextSum[-7]~6\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|NextSum[-7]~6_combout\ = (!\TheRxFsk|Lowpass|Add4~5_sumout\ & (\TheRxFsk|Lowpass|Add4~1_sumout\ & \TheRxFsk|Lowpass|Add4~33_sumout\)) # (\TheRxFsk|Lowpass|Add4~5_sumout\ & ((\TheRxFsk|Lowpass|Add4~33_sumout\) # 
-- (\TheRxFsk|Lowpass|Add4~1_sumout\)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001011100010111000101110001011100010111000101110001011100010111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_Add4~5_sumout\,
	datab => \TheRxFsk|Lowpass|ALT_INV_Add4~1_sumout\,
	datac => \TheRxFsk|Lowpass|ALT_INV_Add4~33_sumout\,
	combout => \TheRxFsk|Lowpass|NextSum[-7]~6_combout\);

-- Location: FF_X30_Y62_N52
\TheRxFsk|Lowpass|Sum[-7]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|NextSum[-7]~6_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Lowpass|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Lowpass|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|Sum[-7]~q\);

-- Location: LABCELL_X31_Y62_N27
\TheRxFsk|Lowpass|Add4~29\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add4~29_sumout\ = SUM(( \TheRxFsk|Lowpass|Sum[-6]~q\ ) + ( \TheRxFsk|Lowpass|MultResult[-6]~5_combout\ ) + ( \TheRxFsk|Lowpass|Add4~34\ ))
-- \TheRxFsk|Lowpass|Add4~30\ = CARRY(( \TheRxFsk|Lowpass|Sum[-6]~q\ ) + ( \TheRxFsk|Lowpass|MultResult[-6]~5_combout\ ) + ( \TheRxFsk|Lowpass|Add4~34\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000101010101010101000000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_MultResult[-6]~5_combout\,
	datac => \TheRxFsk|Lowpass|ALT_INV_Sum[-6]~q\,
	cin => \TheRxFsk|Lowpass|Add4~34\,
	sumout => \TheRxFsk|Lowpass|Add4~29_sumout\,
	cout => \TheRxFsk|Lowpass|Add4~30\);

-- Location: LABCELL_X30_Y62_N48
\TheRxFsk|Lowpass|NextSum[-6]~5\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|NextSum[-6]~5_combout\ = (!\TheRxFsk|Lowpass|Add4~5_sumout\ & (\TheRxFsk|Lowpass|Add4~1_sumout\ & \TheRxFsk|Lowpass|Add4~29_sumout\)) # (\TheRxFsk|Lowpass|Add4~5_sumout\ & ((\TheRxFsk|Lowpass|Add4~29_sumout\) # 
-- (\TheRxFsk|Lowpass|Add4~1_sumout\)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001011100010111000101110001011100010111000101110001011100010111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_Add4~5_sumout\,
	datab => \TheRxFsk|Lowpass|ALT_INV_Add4~1_sumout\,
	datac => \TheRxFsk|Lowpass|ALT_INV_Add4~29_sumout\,
	combout => \TheRxFsk|Lowpass|NextSum[-6]~5_combout\);

-- Location: FF_X30_Y62_N49
\TheRxFsk|Lowpass|Sum[-6]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|NextSum[-6]~5_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Lowpass|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Lowpass|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|Sum[-6]~q\);

-- Location: LABCELL_X31_Y62_N30
\TheRxFsk|Lowpass|Add4~25\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add4~25_sumout\ = SUM(( \TheRxFsk|Lowpass|Sum[-5]~q\ ) + ( \TheRxFsk|Lowpass|MultResult[-5]~4_combout\ ) + ( \TheRxFsk|Lowpass|Add4~30\ ))
-- \TheRxFsk|Lowpass|Add4~26\ = CARRY(( \TheRxFsk|Lowpass|Sum[-5]~q\ ) + ( \TheRxFsk|Lowpass|MultResult[-5]~4_combout\ ) + ( \TheRxFsk|Lowpass|Add4~30\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000110011001100110000000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Lowpass|ALT_INV_MultResult[-5]~4_combout\,
	datac => \TheRxFsk|Lowpass|ALT_INV_Sum[-5]~q\,
	cin => \TheRxFsk|Lowpass|Add4~30\,
	sumout => \TheRxFsk|Lowpass|Add4~25_sumout\,
	cout => \TheRxFsk|Lowpass|Add4~26\);

-- Location: LABCELL_X30_Y62_N21
\TheRxFsk|Lowpass|NextSum[-5]~4\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|NextSum[-5]~4_combout\ = ( \TheRxFsk|Lowpass|Add4~25_sumout\ & ( (\TheRxFsk|Lowpass|Add4~1_sumout\) # (\TheRxFsk|Lowpass|Add4~5_sumout\) ) ) # ( !\TheRxFsk|Lowpass|Add4~25_sumout\ & ( (\TheRxFsk|Lowpass|Add4~5_sumout\ & 
-- \TheRxFsk|Lowpass|Add4~1_sumout\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000100010001000100010001000101110111011101110111011101110111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_Add4~5_sumout\,
	datab => \TheRxFsk|Lowpass|ALT_INV_Add4~1_sumout\,
	dataf => \TheRxFsk|Lowpass|ALT_INV_Add4~25_sumout\,
	combout => \TheRxFsk|Lowpass|NextSum[-5]~4_combout\);

-- Location: FF_X30_Y62_N22
\TheRxFsk|Lowpass|Sum[-5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|NextSum[-5]~4_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Lowpass|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Lowpass|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|Sum[-5]~q\);

-- Location: LABCELL_X31_Y62_N33
\TheRxFsk|Lowpass|Add4~21\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add4~21_sumout\ = SUM(( \TheRxFsk|Lowpass|Sum[-4]~q\ ) + ( \TheRxFsk|Lowpass|MultResult[-4]~3_combout\ ) + ( \TheRxFsk|Lowpass|Add4~26\ ))
-- \TheRxFsk|Lowpass|Add4~22\ = CARRY(( \TheRxFsk|Lowpass|Sum[-4]~q\ ) + ( \TheRxFsk|Lowpass|MultResult[-4]~3_combout\ ) + ( \TheRxFsk|Lowpass|Add4~26\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111110000000000000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Lowpass|ALT_INV_Sum[-4]~q\,
	dataf => \TheRxFsk|Lowpass|ALT_INV_MultResult[-4]~3_combout\,
	cin => \TheRxFsk|Lowpass|Add4~26\,
	sumout => \TheRxFsk|Lowpass|Add4~21_sumout\,
	cout => \TheRxFsk|Lowpass|Add4~22\);

-- Location: LABCELL_X30_Y62_N18
\TheRxFsk|Lowpass|NextSum[-4]~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|NextSum[-4]~3_combout\ = (!\TheRxFsk|Lowpass|Add4~5_sumout\ & (\TheRxFsk|Lowpass|Add4~1_sumout\ & \TheRxFsk|Lowpass|Add4~21_sumout\)) # (\TheRxFsk|Lowpass|Add4~5_sumout\ & ((\TheRxFsk|Lowpass|Add4~21_sumout\) # 
-- (\TheRxFsk|Lowpass|Add4~1_sumout\)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001011100010111000101110001011100010111000101110001011100010111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_Add4~5_sumout\,
	datab => \TheRxFsk|Lowpass|ALT_INV_Add4~1_sumout\,
	datac => \TheRxFsk|Lowpass|ALT_INV_Add4~21_sumout\,
	combout => \TheRxFsk|Lowpass|NextSum[-4]~3_combout\);

-- Location: FF_X30_Y62_N19
\TheRxFsk|Lowpass|Sum[-4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|NextSum[-4]~3_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Lowpass|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Lowpass|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|Sum[-4]~q\);

-- Location: LABCELL_X31_Y62_N36
\TheRxFsk|Lowpass|Add4~17\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add4~17_sumout\ = SUM(( \TheRxFsk|Lowpass|Sum[-3]~q\ ) + ( \TheRxFsk|Lowpass|MultResult[-3]~2_combout\ ) + ( \TheRxFsk|Lowpass|Add4~22\ ))
-- \TheRxFsk|Lowpass|Add4~18\ = CARRY(( \TheRxFsk|Lowpass|Sum[-3]~q\ ) + ( \TheRxFsk|Lowpass|MultResult[-3]~2_combout\ ) + ( \TheRxFsk|Lowpass|Add4~22\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000101010101010101000000000000000000011001100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_MultResult[-3]~2_combout\,
	datab => \TheRxFsk|Lowpass|ALT_INV_Sum[-3]~q\,
	cin => \TheRxFsk|Lowpass|Add4~22\,
	sumout => \TheRxFsk|Lowpass|Add4~17_sumout\,
	cout => \TheRxFsk|Lowpass|Add4~18\);

-- Location: LABCELL_X30_Y62_N3
\TheRxFsk|Lowpass|NextSum[-3]~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|NextSum[-3]~2_combout\ = (!\TheRxFsk|Lowpass|Add4~5_sumout\ & (\TheRxFsk|Lowpass|Add4~1_sumout\ & \TheRxFsk|Lowpass|Add4~17_sumout\)) # (\TheRxFsk|Lowpass|Add4~5_sumout\ & ((\TheRxFsk|Lowpass|Add4~17_sumout\) # 
-- (\TheRxFsk|Lowpass|Add4~1_sumout\)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001011100010111000101110001011100010111000101110001011100010111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_Add4~5_sumout\,
	datab => \TheRxFsk|Lowpass|ALT_INV_Add4~1_sumout\,
	datac => \TheRxFsk|Lowpass|ALT_INV_Add4~17_sumout\,
	combout => \TheRxFsk|Lowpass|NextSum[-3]~2_combout\);

-- Location: FF_X30_Y62_N4
\TheRxFsk|Lowpass|Sum[-3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|NextSum[-3]~2_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Lowpass|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Lowpass|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|Sum[-3]~q\);

-- Location: LABCELL_X31_Y62_N39
\TheRxFsk|Lowpass|Add4~13\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add4~13_sumout\ = SUM(( \TheRxFsk|Lowpass|Sum[-2]~q\ ) + ( \TheRxFsk|Lowpass|MultResult[-2]~1_combout\ ) + ( \TheRxFsk|Lowpass|Add4~18\ ))
-- \TheRxFsk|Lowpass|Add4~14\ = CARRY(( \TheRxFsk|Lowpass|Sum[-2]~q\ ) + ( \TheRxFsk|Lowpass|MultResult[-2]~1_combout\ ) + ( \TheRxFsk|Lowpass|Add4~18\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000111111110000000000000000000000000000111100001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Lowpass|ALT_INV_Sum[-2]~q\,
	dataf => \TheRxFsk|Lowpass|ALT_INV_MultResult[-2]~1_combout\,
	cin => \TheRxFsk|Lowpass|Add4~18\,
	sumout => \TheRxFsk|Lowpass|Add4~13_sumout\,
	cout => \TheRxFsk|Lowpass|Add4~14\);

-- Location: LABCELL_X30_Y62_N0
\TheRxFsk|Lowpass|NextSum[-2]~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|NextSum[-2]~1_combout\ = (!\TheRxFsk|Lowpass|Add4~5_sumout\ & (\TheRxFsk|Lowpass|Add4~1_sumout\ & \TheRxFsk|Lowpass|Add4~13_sumout\)) # (\TheRxFsk|Lowpass|Add4~5_sumout\ & ((\TheRxFsk|Lowpass|Add4~13_sumout\) # 
-- (\TheRxFsk|Lowpass|Add4~1_sumout\)))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001011100010111000101110001011100010111000101110001011100010111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_Add4~5_sumout\,
	datab => \TheRxFsk|Lowpass|ALT_INV_Add4~1_sumout\,
	datac => \TheRxFsk|Lowpass|ALT_INV_Add4~13_sumout\,
	combout => \TheRxFsk|Lowpass|NextSum[-2]~1_combout\);

-- Location: FF_X30_Y62_N1
\TheRxFsk|Lowpass|Sum[-2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|NextSum[-2]~1_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Lowpass|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Lowpass|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|Sum[-2]~q\);

-- Location: LABCELL_X31_Y62_N42
\TheRxFsk|Lowpass|Add4~9\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add4~9_sumout\ = SUM(( \TheRxFsk|Lowpass|MultResult[-1]~0_combout\ ) + ( \TheRxFsk|Lowpass|Sum[-1]~q\ ) + ( \TheRxFsk|Lowpass|Add4~14\ ))
-- \TheRxFsk|Lowpass|Add4~10\ = CARRY(( \TheRxFsk|Lowpass|MultResult[-1]~0_combout\ ) + ( \TheRxFsk|Lowpass|Sum[-1]~q\ ) + ( \TheRxFsk|Lowpass|Add4~14\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000110011001100110000000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Lowpass|ALT_INV_Sum[-1]~q\,
	datad => \TheRxFsk|Lowpass|ALT_INV_MultResult[-1]~0_combout\,
	cin => \TheRxFsk|Lowpass|Add4~14\,
	sumout => \TheRxFsk|Lowpass|Add4~9_sumout\,
	cout => \TheRxFsk|Lowpass|Add4~10\);

-- Location: LABCELL_X30_Y62_N33
\TheRxFsk|Lowpass|NextSum[-1]~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|NextSum[-1]~0_combout\ = ( \TheRxFsk|Lowpass|Add4~9_sumout\ & ( \TheRxFsk|Lowpass|Add4~5_sumout\ ) ) # ( !\TheRxFsk|Lowpass|Add4~9_sumout\ & ( \TheRxFsk|Lowpass|Add4~5_sumout\ & ( \TheRxFsk|Lowpass|Add4~1_sumout\ ) ) ) # ( 
-- \TheRxFsk|Lowpass|Add4~9_sumout\ & ( !\TheRxFsk|Lowpass|Add4~5_sumout\ & ( \TheRxFsk|Lowpass|Add4~1_sumout\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000011110000111100001111000011111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheRxFsk|Lowpass|ALT_INV_Add4~1_sumout\,
	datae => \TheRxFsk|Lowpass|ALT_INV_Add4~9_sumout\,
	dataf => \TheRxFsk|Lowpass|ALT_INV_Add4~5_sumout\,
	combout => \TheRxFsk|Lowpass|NextSum[-1]~0_combout\);

-- Location: FF_X30_Y62_N34
\TheRxFsk|Lowpass|Sum[-1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|NextSum[-1]~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Lowpass|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Lowpass|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|Sum[-1]~q\);

-- Location: LABCELL_X31_Y62_N48
\TheRxFsk|Lowpass|Add4~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add4~1_sumout\ = SUM(( \TheRxFsk|Lowpass|Sum\(0) ) + ( !\TheRxFsk|Lowpass|MultResultDelayed\(0) ) + ( \TheRxFsk|Lowpass|Add4~6\ ))

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000001100110011001100000000000000000000000011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Lowpass|ALT_INV_MultResultDelayed\(0),
	datad => \TheRxFsk|Lowpass|ALT_INV_Sum\(0),
	cin => \TheRxFsk|Lowpass|Add4~6\,
	sumout => \TheRxFsk|Lowpass|Add4~1_sumout\);

-- Location: LABCELL_X30_Y62_N36
\TheRxFsk|Lowpass|Add4~1_wirecell\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Add4~1_wirecell_combout\ = ( !\TheRxFsk|Lowpass|Add4~1_sumout\ )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111111111111111000000000000000011111111111111110000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datae => \TheRxFsk|Lowpass|ALT_INV_Add4~1_sumout\,
	combout => \TheRxFsk|Lowpass|Add4~1_wirecell_combout\);

-- Location: FF_X30_Y62_N37
\TheRxFsk|Lowpass|Sum[0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|Add4~1_wirecell_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sclr => \TheRxFsk|Lowpass|ALT_INV_R.SelSumUp~q\,
	ena => \TheRxFsk|Lowpass|R.EnableSumUp~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|Sum\(0));

-- Location: LABCELL_X31_Y60_N24
\TheRxFsk|Lowpass|Selector8~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|Lowpass|Selector8~0_combout\ = ( \TheRxFsk|Lowpass|R.SumState.SumWait2~DUPLICATE_q\ ) # ( !\TheRxFsk|Lowpass|R.SumState.SumWait2~DUPLICATE_q\ & ( (!\TheRxFsk|Lowpass|R.SumState.SumValid~q\ & \TheRxFsk|Lowpass|R.ValWet~q\) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011001100000000001100110011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheRxFsk|Lowpass|ALT_INV_R.SumState.SumValid~q\,
	datad => \TheRxFsk|Lowpass|ALT_INV_R.ValWet~q\,
	dataf => \TheRxFsk|Lowpass|ALT_INV_R.SumState.SumWait2~DUPLICATE_q\,
	combout => \TheRxFsk|Lowpass|Selector8~0_combout\);

-- Location: FF_X31_Y60_N25
\TheRxFsk|Lowpass|R.ValWet\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|Lowpass|Selector8~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|Lowpass|R.ValWet~q\);

-- Location: LABCELL_X31_Y60_N27
\TheRxFsk|oD~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheRxFsk|oD~0_combout\ = ( \TheRxFsk|Lowpass|R.ValWet~q\ & ( !\TheRxFsk|Lowpass|Sum\(0) ) ) # ( !\TheRxFsk|Lowpass|R.ValWet~q\ & ( \TheRxFsk|oD~q\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011111111000000001111111110101010101010101010101010101010",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheRxFsk|Lowpass|ALT_INV_Sum\(0),
	datad => \TheRxFsk|ALT_INV_oD~q\,
	dataf => \TheRxFsk|Lowpass|ALT_INV_R.ValWet~q\,
	combout => \TheRxFsk|oD~0_combout\);

-- Location: FF_X31_Y60_N28
\TheRxFsk|oD\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \iClk~inputCLKENA0_outclk\,
	d => \TheRxFsk|oD~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheRxFsk|oD~q\);

-- Location: FF_X13_Y63_N50
\TheParToI2s|BclkCtr[3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \TheParToI2s|Selector6~2_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheParToI2s|BclkCtr\(3));

-- Location: LABCELL_X13_Y64_N42
\TheParToI2s|Selector0~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheParToI2s|Selector0~0_combout\ = ( \TheParToI2s|State.WaitingValL~q\ & ( \TheParToI2s|State.SendingR~q\ & ( !\TheParToI2s|NextState~6_combout\ ) ) ) # ( !\TheParToI2s|State.WaitingValL~q\ & ( \TheParToI2s|State.SendingR~q\ & ( 
-- (!\TheParToI2s|NextState~6_combout\ & \TheI2sToPar|ValL~q\) ) ) ) # ( \TheParToI2s|State.WaitingValL~q\ & ( !\TheParToI2s|State.SendingR~q\ ) ) # ( !\TheParToI2s|State.WaitingValL~q\ & ( !\TheParToI2s|State.SendingR~q\ & ( \TheI2sToPar|ValL~q\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111111111111111111100001100000011001100110011001100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datab => \TheParToI2s|ALT_INV_NextState~6_combout\,
	datac => \TheI2sToPar|ALT_INV_ValL~q\,
	datae => \TheParToI2s|ALT_INV_State.WaitingValL~q\,
	dataf => \TheParToI2s|ALT_INV_State.SendingR~q\,
	combout => \TheParToI2s|Selector0~0_combout\);

-- Location: FF_X13_Y64_N43
\TheParToI2s|State.WaitingValL\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \TheParToI2s|Selector0~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheParToI2s|State.WaitingValL~q\);

-- Location: LABCELL_X13_Y63_N30
\TheParToI2s|Selector1~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheParToI2s|Selector1~0_combout\ = ( \TheI2sToPar|ValL~q\ & ( (!\TheParToI2s|State.WaitingValL~q\) # ((\TheParToI2s|State.SyncingToBclk~q\ & ((!\TheI2sToPar|BclkDlyd~q\) # (\GenClks|BMclk~q\)))) ) ) # ( !\TheI2sToPar|ValL~q\ & ( 
-- (\TheParToI2s|State.SyncingToBclk~q\ & ((!\TheI2sToPar|BclkDlyd~q\) # (\GenClks|BMclk~q\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000010111011000000001011101111110000111110111111000011111011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheI2sToPar|ALT_INV_BclkDlyd~q\,
	datab => \GenClks|ALT_INV_BMclk~q\,
	datac => \TheParToI2s|ALT_INV_State.WaitingValL~q\,
	datad => \TheParToI2s|ALT_INV_State.SyncingToBclk~q\,
	dataf => \TheI2sToPar|ALT_INV_ValL~q\,
	combout => \TheParToI2s|Selector1~0_combout\);

-- Location: FF_X13_Y63_N31
\TheParToI2s|State.SyncingToBclk\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \TheParToI2s|Selector1~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheParToI2s|State.SyncingToBclk~q\);

-- Location: LABCELL_X13_Y63_N33
\TheParToI2s|State.FirstBitEmptyL~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheParToI2s|State.FirstBitEmptyL~0_combout\ = ( \TheParToI2s|State.SyncingToBclk~q\ & ( ((\TheI2sToPar|BclkDlyd~q\ & !\GenClks|BMclk~q\)) # (\TheParToI2s|State.FirstBitEmptyL~q\) ) ) # ( !\TheParToI2s|State.SyncingToBclk~q\ & ( 
-- (\TheParToI2s|State.FirstBitEmptyL~q\ & ((!\TheI2sToPar|BclkDlyd~q\) # (\GenClks|BMclk~q\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000010111011000000001011101101000100111111110100010011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheI2sToPar|ALT_INV_BclkDlyd~q\,
	datab => \GenClks|ALT_INV_BMclk~q\,
	datad => \TheParToI2s|ALT_INV_State.FirstBitEmptyL~q\,
	dataf => \TheParToI2s|ALT_INV_State.SyncingToBclk~q\,
	combout => \TheParToI2s|State.FirstBitEmptyL~0_combout\);

-- Location: FF_X13_Y63_N35
\TheParToI2s|State.FirstBitEmptyL\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \TheParToI2s|State.FirstBitEmptyL~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheParToI2s|State.FirstBitEmptyL~q\);

-- Location: LABCELL_X13_Y64_N51
\TheParToI2s|Selector3~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheParToI2s|Selector3~0_combout\ = ( \TheParToI2s|State.SendingL~q\ & ( \TheParToI2s|NextState~6_combout\ & ( (\TheI2sToPar|BclkDlyd~q\ & (\TheParToI2s|State.FirstBitEmptyL~q\ & !\GenClks|BMclk~q\)) ) ) ) # ( !\TheParToI2s|State.SendingL~q\ & ( 
-- \TheParToI2s|NextState~6_combout\ & ( (\TheI2sToPar|BclkDlyd~q\ & (\TheParToI2s|State.FirstBitEmptyL~q\ & !\GenClks|BMclk~q\)) ) ) ) # ( \TheParToI2s|State.SendingL~q\ & ( !\TheParToI2s|NextState~6_combout\ ) ) # ( !\TheParToI2s|State.SendingL~q\ & ( 
-- !\TheParToI2s|NextState~6_combout\ & ( (\TheI2sToPar|BclkDlyd~q\ & (\TheParToI2s|State.FirstBitEmptyL~q\ & !\GenClks|BMclk~q\)) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001000000010000111111111111111100010000000100000001000000010000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheI2sToPar|ALT_INV_BclkDlyd~q\,
	datab => \TheParToI2s|ALT_INV_State.FirstBitEmptyL~q\,
	datac => \GenClks|ALT_INV_BMclk~q\,
	datae => \TheParToI2s|ALT_INV_State.SendingL~q\,
	dataf => \TheParToI2s|ALT_INV_NextState~6_combout\,
	combout => \TheParToI2s|Selector3~0_combout\);

-- Location: FF_X13_Y64_N52
\TheParToI2s|State.SendingL\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \TheParToI2s|Selector3~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheParToI2s|State.SendingL~q\);

-- Location: LABCELL_X13_Y64_N57
\TheParToI2s|Selector4~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheParToI2s|Selector4~0_combout\ = ( \TheParToI2s|State.FirstBitEmptyR~q\ & ( \TheParToI2s|State.SendingL~q\ & ( (!\TheI2sToPar|BclkDlyd~q\) # ((\GenClks|BMclk~q\) # (\TheParToI2s|NextState~6_combout\)) ) ) ) # ( !\TheParToI2s|State.FirstBitEmptyR~q\ & ( 
-- \TheParToI2s|State.SendingL~q\ & ( \TheParToI2s|NextState~6_combout\ ) ) ) # ( \TheParToI2s|State.FirstBitEmptyR~q\ & ( !\TheParToI2s|State.SendingL~q\ & ( (!\TheI2sToPar|BclkDlyd~q\) # (\GenClks|BMclk~q\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000101011111010111100110011001100111011111110111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheI2sToPar|ALT_INV_BclkDlyd~q\,
	datab => \TheParToI2s|ALT_INV_NextState~6_combout\,
	datac => \GenClks|ALT_INV_BMclk~q\,
	datae => \TheParToI2s|ALT_INV_State.FirstBitEmptyR~q\,
	dataf => \TheParToI2s|ALT_INV_State.SendingL~q\,
	combout => \TheParToI2s|Selector4~0_combout\);

-- Location: FF_X13_Y64_N58
\TheParToI2s|State.FirstBitEmptyR\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \TheParToI2s|Selector4~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheParToI2s|State.FirstBitEmptyR~q\);

-- Location: LABCELL_X13_Y63_N27
\TheParToI2s|Selector8~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheParToI2s|Selector8~0_combout\ = ( \TheParToI2s|State.FirstBitEmptyL~q\ & ( ((\TheI2sToPar|BclkDlyd~q\ & !\GenClks|BMclk~q\)) # (\TheParToI2s|BclkCtr\(1)) ) ) # ( !\TheParToI2s|State.FirstBitEmptyL~q\ & ( (\TheParToI2s|State.FirstBitEmptyR~q\ & 
-- (((\TheI2sToPar|BclkDlyd~q\ & !\GenClks|BMclk~q\)) # (\TheParToI2s|BclkCtr\(1)))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000011100000011000001110000001101110111001100110111011100110011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheI2sToPar|ALT_INV_BclkDlyd~q\,
	datab => \TheParToI2s|ALT_INV_BclkCtr\(1),
	datac => \TheParToI2s|ALT_INV_State.FirstBitEmptyR~q\,
	datad => \GenClks|ALT_INV_BMclk~q\,
	dataf => \TheParToI2s|ALT_INV_State.FirstBitEmptyL~q\,
	combout => \TheParToI2s|Selector8~0_combout\);

-- Location: FF_X13_Y63_N32
\TheParToI2s|State.SyncingToBclk~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \TheParToI2s|Selector1~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheParToI2s|State.SyncingToBclk~DUPLICATE_q\);

-- Location: LABCELL_X13_Y63_N21
\TheParToI2s|NextBclkCtr~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheParToI2s|NextBclkCtr~0_combout\ = (!\TheParToI2s|State.SyncingToBclk~DUPLICATE_q\ & \TheParToI2s|State.WaitingValL~q\)

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011110000000000001111000000000000111100000000000011110000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheParToI2s|ALT_INV_State.SyncingToBclk~DUPLICATE_q\,
	datad => \TheParToI2s|ALT_INV_State.WaitingValL~q\,
	combout => \TheParToI2s|NextBclkCtr~0_combout\);

-- Location: LABCELL_X13_Y63_N3
\TheParToI2s|Selector7~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheParToI2s|Selector7~0_combout\ = ( \GenClks|BMclk~q\ & ( (\TheParToI2s|BclkCtr\(2) & ((\TheParToI2s|State.FirstBitEmptyR~q\) # (\TheParToI2s|State.FirstBitEmptyL~q\))) ) ) # ( !\GenClks|BMclk~q\ & ( (!\TheParToI2s|State.FirstBitEmptyL~q\ & 
-- (\TheParToI2s|State.FirstBitEmptyR~q\ & ((\TheI2sToPar|BclkDlyd~q\) # (\TheParToI2s|BclkCtr\(2))))) # (\TheParToI2s|State.FirstBitEmptyL~q\ & (((\TheI2sToPar|BclkDlyd~q\)) # (\TheParToI2s|BclkCtr\(2)))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001001101011111000100110101111100010011000100110001001100010011",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheParToI2s|ALT_INV_State.FirstBitEmptyL~q\,
	datab => \TheParToI2s|ALT_INV_BclkCtr\(2),
	datac => \TheParToI2s|ALT_INV_State.FirstBitEmptyR~q\,
	datad => \TheI2sToPar|ALT_INV_BclkDlyd~q\,
	dataf => \GenClks|ALT_INV_BMclk~q\,
	combout => \TheParToI2s|Selector7~0_combout\);

-- Location: LABCELL_X13_Y63_N18
\TheParToI2s|Selector9~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheParToI2s|Selector9~0_combout\ = ( \TheParToI2s|State.FirstBitEmptyR~q\ & ( ((\TheI2sToPar|BclkDlyd~q\ & !\GenClks|BMclk~q\)) # (\TheParToI2s|BclkCtr\(0)) ) ) # ( !\TheParToI2s|State.FirstBitEmptyR~q\ & ( (\TheParToI2s|State.FirstBitEmptyL~q\ & 
-- (((\TheI2sToPar|BclkDlyd~q\ & !\GenClks|BMclk~q\)) # (\TheParToI2s|BclkCtr\(0)))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010000001111000001000000111101000100111111110100010011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheI2sToPar|ALT_INV_BclkDlyd~q\,
	datab => \GenClks|ALT_INV_BMclk~q\,
	datac => \TheParToI2s|ALT_INV_State.FirstBitEmptyL~q\,
	datad => \TheParToI2s|ALT_INV_BclkCtr\(0),
	dataf => \TheParToI2s|ALT_INV_State.FirstBitEmptyR~q\,
	combout => \TheParToI2s|Selector9~0_combout\);

-- Location: LABCELL_X13_Y63_N51
\TheParToI2s|Selector9~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheParToI2s|Selector9~1_combout\ = ( \TheParToI2s|Selector9~0_combout\ ) # ( !\TheParToI2s|Selector9~0_combout\ & ( (!\TheParToI2s|BclkCtr\(0) & (\TheParToI2s|Selector10~0_combout\ & ((\TheParToI2s|NextBclkCtr~1_combout\)))) # (\TheParToI2s|BclkCtr\(0) & 
-- ((!\TheParToI2s|NextBclkCtr~0_combout\) # ((\TheParToI2s|Selector10~0_combout\ & !\TheParToI2s|NextBclkCtr~1_combout\)))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010111011100000001011101110011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheParToI2s|ALT_INV_Selector10~0_combout\,
	datab => \TheParToI2s|ALT_INV_NextBclkCtr~0_combout\,
	datac => \TheParToI2s|ALT_INV_NextBclkCtr~1_combout\,
	datad => \TheParToI2s|ALT_INV_BclkCtr\(0),
	dataf => \TheParToI2s|ALT_INV_Selector9~0_combout\,
	combout => \TheParToI2s|Selector9~1_combout\);

-- Location: FF_X13_Y63_N52
\TheParToI2s|BclkCtr[0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \TheParToI2s|Selector9~1_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheParToI2s|BclkCtr\(0));

-- Location: LABCELL_X13_Y63_N24
\TheParToI2s|Add0~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheParToI2s|Add0~0_combout\ = ( !\TheParToI2s|BclkCtr\(1) & ( !\TheParToI2s|BclkCtr\(0) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "1111000011110000111100001111000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheParToI2s|ALT_INV_BclkCtr\(0),
	dataf => \TheParToI2s|ALT_INV_BclkCtr\(1),
	combout => \TheParToI2s|Add0~0_combout\);

-- Location: LABCELL_X13_Y63_N12
\TheParToI2s|Selector7~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheParToI2s|Selector7~1_combout\ = ( \TheParToI2s|BclkCtr\(2) & ( \TheParToI2s|Add0~0_combout\ & ( (!\TheParToI2s|NextBclkCtr~0_combout\) # (((\TheParToI2s|Selector10~0_combout\ & !\TheParToI2s|NextBclkCtr~1_combout\)) # 
-- (\TheParToI2s|Selector7~0_combout\)) ) ) ) # ( !\TheParToI2s|BclkCtr\(2) & ( \TheParToI2s|Add0~0_combout\ & ( ((\TheParToI2s|Selector10~0_combout\ & \TheParToI2s|NextBclkCtr~1_combout\)) # (\TheParToI2s|Selector7~0_combout\) ) ) ) # ( 
-- \TheParToI2s|BclkCtr\(2) & ( !\TheParToI2s|Add0~0_combout\ & ( ((!\TheParToI2s|NextBclkCtr~0_combout\) # (\TheParToI2s|Selector7~0_combout\)) # (\TheParToI2s|Selector10~0_combout\) ) ) ) # ( !\TheParToI2s|BclkCtr\(2) & ( !\TheParToI2s|Add0~0_combout\ & ( 
-- \TheParToI2s|Selector7~0_combout\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111110111111101111100001111010111111101111111001111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheParToI2s|ALT_INV_Selector10~0_combout\,
	datab => \TheParToI2s|ALT_INV_NextBclkCtr~0_combout\,
	datac => \TheParToI2s|ALT_INV_Selector7~0_combout\,
	datad => \TheParToI2s|ALT_INV_NextBclkCtr~1_combout\,
	datae => \TheParToI2s|ALT_INV_BclkCtr\(2),
	dataf => \TheParToI2s|ALT_INV_Add0~0_combout\,
	combout => \TheParToI2s|Selector7~1_combout\);

-- Location: FF_X13_Y63_N14
\TheParToI2s|BclkCtr[2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \TheParToI2s|Selector7~1_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheParToI2s|BclkCtr\(2));

-- Location: LABCELL_X13_Y63_N39
\TheParToI2s|NextBclkCtr~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheParToI2s|NextBclkCtr~1_combout\ = ( \TheParToI2s|BclkCtr[3]~DUPLICATE_q\ & ( \TheParToI2s|BclkCtr\(1) & ( (\TheI2sToPar|BclkDlyd~q\ & !\GenClks|BMclk~q\) ) ) ) # ( !\TheParToI2s|BclkCtr[3]~DUPLICATE_q\ & ( \TheParToI2s|BclkCtr\(1) & ( 
-- (\TheI2sToPar|BclkDlyd~q\ & !\GenClks|BMclk~q\) ) ) ) # ( \TheParToI2s|BclkCtr[3]~DUPLICATE_q\ & ( !\TheParToI2s|BclkCtr\(1) & ( (\TheI2sToPar|BclkDlyd~q\ & !\GenClks|BMclk~q\) ) ) ) # ( !\TheParToI2s|BclkCtr[3]~DUPLICATE_q\ & ( !\TheParToI2s|BclkCtr\(1) 
-- & ( (\TheI2sToPar|BclkDlyd~q\ & (!\GenClks|BMclk~q\ & ((\TheParToI2s|BclkCtr\(0)) # (\TheParToI2s|BclkCtr\(2))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010001000100010001000100010001000100010001000100010001000100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheI2sToPar|ALT_INV_BclkDlyd~q\,
	datab => \GenClks|ALT_INV_BMclk~q\,
	datac => \TheParToI2s|ALT_INV_BclkCtr\(2),
	datad => \TheParToI2s|ALT_INV_BclkCtr\(0),
	datae => \TheParToI2s|ALT_INV_BclkCtr[3]~DUPLICATE_q\,
	dataf => \TheParToI2s|ALT_INV_BclkCtr\(1),
	combout => \TheParToI2s|NextBclkCtr~1_combout\);

-- Location: LABCELL_X13_Y63_N45
\TheParToI2s|Selector8~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheParToI2s|Selector8~1_combout\ = ( \TheParToI2s|BclkCtr\(1) & ( \TheParToI2s|BclkCtr\(0) & ( ((!\TheParToI2s|NextBclkCtr~0_combout\) # (\TheParToI2s|Selector10~0_combout\)) # (\TheParToI2s|Selector8~0_combout\) ) ) ) # ( !\TheParToI2s|BclkCtr\(1) & ( 
-- \TheParToI2s|BclkCtr\(0) & ( \TheParToI2s|Selector8~0_combout\ ) ) ) # ( \TheParToI2s|BclkCtr\(1) & ( !\TheParToI2s|BclkCtr\(0) & ( ((!\TheParToI2s|NextBclkCtr~0_combout\) # ((!\TheParToI2s|NextBclkCtr~1_combout\ & \TheParToI2s|Selector10~0_combout\))) # 
-- (\TheParToI2s|Selector8~0_combout\) ) ) ) # ( !\TheParToI2s|BclkCtr\(1) & ( !\TheParToI2s|BclkCtr\(0) & ( ((\TheParToI2s|NextBclkCtr~1_combout\ & \TheParToI2s|Selector10~0_combout\)) # (\TheParToI2s|Selector8~0_combout\) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010101110111111101011111110101010101010101011111010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheParToI2s|ALT_INV_Selector8~0_combout\,
	datab => \TheParToI2s|ALT_INV_NextBclkCtr~1_combout\,
	datac => \TheParToI2s|ALT_INV_NextBclkCtr~0_combout\,
	datad => \TheParToI2s|ALT_INV_Selector10~0_combout\,
	datae => \TheParToI2s|ALT_INV_BclkCtr\(1),
	dataf => \TheParToI2s|ALT_INV_BclkCtr\(0),
	combout => \TheParToI2s|Selector8~1_combout\);

-- Location: FF_X13_Y63_N46
\TheParToI2s|BclkCtr[1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \TheParToI2s|Selector8~1_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheParToI2s|BclkCtr\(1));

-- Location: LABCELL_X13_Y63_N9
\TheParToI2s|NextState~6\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheParToI2s|NextState~6_combout\ = ( \TheI2sToPar|BclkDlyd~q\ & ( !\TheParToI2s|BclkCtr\(2) & ( (!\TheParToI2s|BclkCtr\(3) & (!\GenClks|BMclk~q\ & (!\TheParToI2s|BclkCtr\(1) & !\TheParToI2s|BclkCtr\(0)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000100000000000000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheParToI2s|ALT_INV_BclkCtr\(3),
	datab => \GenClks|ALT_INV_BMclk~q\,
	datac => \TheParToI2s|ALT_INV_BclkCtr\(1),
	datad => \TheParToI2s|ALT_INV_BclkCtr\(0),
	datae => \TheI2sToPar|ALT_INV_BclkDlyd~q\,
	dataf => \TheParToI2s|ALT_INV_BclkCtr\(2),
	combout => \TheParToI2s|NextState~6_combout\);

-- Location: LABCELL_X13_Y64_N21
\TheParToI2s|Selector5~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheParToI2s|Selector5~0_combout\ = ( \TheParToI2s|State.SendingR~q\ & ( \TheParToI2s|State.FirstBitEmptyR~q\ & ( (!\TheParToI2s|NextState~6_combout\) # ((\TheI2sToPar|BclkDlyd~q\ & !\GenClks|BMclk~q\)) ) ) ) # ( !\TheParToI2s|State.SendingR~q\ & ( 
-- \TheParToI2s|State.FirstBitEmptyR~q\ & ( (\TheI2sToPar|BclkDlyd~q\ & !\GenClks|BMclk~q\) ) ) ) # ( \TheParToI2s|State.SendingR~q\ & ( !\TheParToI2s|State.FirstBitEmptyR~q\ & ( !\TheParToI2s|NextState~6_combout\ ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000110011001100110001010000010100001101110011011100",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheI2sToPar|ALT_INV_BclkDlyd~q\,
	datab => \TheParToI2s|ALT_INV_NextState~6_combout\,
	datac => \GenClks|ALT_INV_BMclk~q\,
	datae => \TheParToI2s|ALT_INV_State.SendingR~q\,
	dataf => \TheParToI2s|ALT_INV_State.FirstBitEmptyR~q\,
	combout => \TheParToI2s|Selector5~0_combout\);

-- Location: FF_X13_Y64_N22
\TheParToI2s|State.SendingR\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \TheParToI2s|Selector5~0_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheParToI2s|State.SendingR~q\);

-- Location: LABCELL_X13_Y64_N30
\TheParToI2s|Selector10~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheParToI2s|Selector10~0_combout\ = ( \TheParToI2s|State.SendingL~q\ ) # ( !\TheParToI2s|State.SendingL~q\ & ( \TheParToI2s|State.SendingR~q\ ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000111100001111000011110000111111111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	datac => \TheParToI2s|ALT_INV_State.SendingR~q\,
	dataf => \TheParToI2s|ALT_INV_State.SendingL~q\,
	combout => \TheParToI2s|Selector10~0_combout\);

-- Location: LABCELL_X13_Y63_N54
\TheParToI2s|Selector6~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheParToI2s|Selector6~1_combout\ = ( !\TheParToI2s|BclkCtr\(2) & ( (\TheI2sToPar|BclkDlyd~q\ & (!\GenClks|BMclk~q\ & (!\TheParToI2s|BclkCtr\(0) & !\TheParToI2s|BclkCtr\(1)))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0100000000000000010000000000000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheI2sToPar|ALT_INV_BclkDlyd~q\,
	datab => \GenClks|ALT_INV_BMclk~q\,
	datac => \TheParToI2s|ALT_INV_BclkCtr\(0),
	datad => \TheParToI2s|ALT_INV_BclkCtr\(1),
	dataf => \TheParToI2s|ALT_INV_BclkCtr\(2),
	combout => \TheParToI2s|Selector6~1_combout\);

-- Location: LABCELL_X13_Y63_N57
\TheParToI2s|Selector6~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheParToI2s|Selector6~0_combout\ = ( \TheParToI2s|State.FirstBitEmptyL~q\ & ( ((\TheI2sToPar|BclkDlyd~q\ & !\GenClks|BMclk~q\)) # (\TheParToI2s|BclkCtr[3]~DUPLICATE_q\) ) ) # ( !\TheParToI2s|State.FirstBitEmptyL~q\ & ( 
-- (\TheParToI2s|State.FirstBitEmptyR~q\ & (((\TheI2sToPar|BclkDlyd~q\ & !\GenClks|BMclk~q\)) # (\TheParToI2s|BclkCtr[3]~DUPLICATE_q\))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000010000001111000001000000111101000100111111110100010011111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheI2sToPar|ALT_INV_BclkDlyd~q\,
	datab => \GenClks|ALT_INV_BMclk~q\,
	datac => \TheParToI2s|ALT_INV_State.FirstBitEmptyR~q\,
	datad => \TheParToI2s|ALT_INV_BclkCtr[3]~DUPLICATE_q\,
	dataf => \TheParToI2s|ALT_INV_State.FirstBitEmptyL~q\,
	combout => \TheParToI2s|Selector6~0_combout\);

-- Location: LABCELL_X13_Y63_N48
\TheParToI2s|Selector6~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheParToI2s|Selector6~2_combout\ = ( \TheParToI2s|Selector6~0_combout\ ) # ( !\TheParToI2s|Selector6~0_combout\ & ( (\TheParToI2s|BclkCtr\(3) & ((!\TheParToI2s|NextBclkCtr~0_combout\) # ((\TheParToI2s|Selector10~0_combout\ & 
-- !\TheParToI2s|Selector6~1_combout\)))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000011011100000000001101110011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheParToI2s|ALT_INV_Selector10~0_combout\,
	datab => \TheParToI2s|ALT_INV_NextBclkCtr~0_combout\,
	datac => \TheParToI2s|ALT_INV_Selector6~1_combout\,
	datad => \TheParToI2s|ALT_INV_BclkCtr\(3),
	dataf => \TheParToI2s|ALT_INV_Selector6~0_combout\,
	combout => \TheParToI2s|Selector6~2_combout\);

-- Location: FF_X13_Y63_N49
\TheParToI2s|BclkCtr[3]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \TheParToI2s|Selector6~2_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheParToI2s|BclkCtr[3]~DUPLICATE_q\);

-- Location: FF_X16_Y65_N50
\TheParToI2s|LastValidDL[4]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	asdata => \TheI2sToPar|D\(4),
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \TheI2sToPar|ValL~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheParToI2s|LastValidDL\(4));

-- Location: LABCELL_X16_Y65_N51
\TheParToI2s|LastValidDL[6]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheParToI2s|LastValidDL[6]~feeder_combout\ = ( \TheI2sToPar|D\(6) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \TheI2sToPar|ALT_INV_D\(6),
	combout => \TheParToI2s|LastValidDL[6]~feeder_combout\);

-- Location: FF_X16_Y65_N52
\TheParToI2s|LastValidDL[6]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \TheParToI2s|LastValidDL[6]~feeder_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	ena => \TheI2sToPar|ValL~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheParToI2s|LastValidDL\(6));

-- Location: FF_X16_Y65_N2
\TheParToI2s|LastValidDL[14]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	asdata => \TheI2sToPar|D\(14),
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \TheI2sToPar|ValL~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheParToI2s|LastValidDL\(14));

-- Location: LABCELL_X16_Y65_N6
\TheParToI2s|LastValidDL[12]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheParToI2s|LastValidDL[12]~feeder_combout\ = ( \TheI2sToPar|D\(12) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \TheI2sToPar|ALT_INV_D\(12),
	combout => \TheParToI2s|LastValidDL[12]~feeder_combout\);

-- Location: FF_X16_Y65_N8
\TheParToI2s|LastValidDL[12]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \TheParToI2s|LastValidDL[12]~feeder_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	ena => \TheI2sToPar|ValL~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheParToI2s|LastValidDL\(12));

-- Location: LABCELL_X16_Y65_N0
\TheParToI2s|Mux1~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheParToI2s|Mux1~1_combout\ = ( \TheParToI2s|LastValidDL\(14) & ( \TheParToI2s|LastValidDL\(12) & ( ((!\TheParToI2s|BclkCtr\(1) & (\TheParToI2s|LastValidDL\(4))) # (\TheParToI2s|BclkCtr\(1) & ((\TheParToI2s|LastValidDL\(6))))) # 
-- (\TheParToI2s|BclkCtr[3]~DUPLICATE_q\) ) ) ) # ( !\TheParToI2s|LastValidDL\(14) & ( \TheParToI2s|LastValidDL\(12) & ( (!\TheParToI2s|BclkCtr[3]~DUPLICATE_q\ & ((!\TheParToI2s|BclkCtr\(1) & (\TheParToI2s|LastValidDL\(4))) # (\TheParToI2s|BclkCtr\(1) & 
-- ((\TheParToI2s|LastValidDL\(6)))))) # (\TheParToI2s|BclkCtr[3]~DUPLICATE_q\ & (!\TheParToI2s|BclkCtr\(1))) ) ) ) # ( \TheParToI2s|LastValidDL\(14) & ( !\TheParToI2s|LastValidDL\(12) & ( (!\TheParToI2s|BclkCtr[3]~DUPLICATE_q\ & ((!\TheParToI2s|BclkCtr\(1) 
-- & (\TheParToI2s|LastValidDL\(4))) # (\TheParToI2s|BclkCtr\(1) & ((\TheParToI2s|LastValidDL\(6)))))) # (\TheParToI2s|BclkCtr[3]~DUPLICATE_q\ & (\TheParToI2s|BclkCtr\(1))) ) ) ) # ( !\TheParToI2s|LastValidDL\(14) & ( !\TheParToI2s|LastValidDL\(12) & ( 
-- (!\TheParToI2s|BclkCtr[3]~DUPLICATE_q\ & ((!\TheParToI2s|BclkCtr\(1) & (\TheParToI2s|LastValidDL\(4))) # (\TheParToI2s|BclkCtr\(1) & ((\TheParToI2s|LastValidDL\(6)))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000100000101010000110010011101101001100011011100101110101111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheParToI2s|ALT_INV_BclkCtr[3]~DUPLICATE_q\,
	datab => \TheParToI2s|ALT_INV_BclkCtr\(1),
	datac => \TheParToI2s|ALT_INV_LastValidDL\(4),
	datad => \TheParToI2s|ALT_INV_LastValidDL\(6),
	datae => \TheParToI2s|ALT_INV_LastValidDL\(14),
	dataf => \TheParToI2s|ALT_INV_LastValidDL\(12),
	combout => \TheParToI2s|Mux1~1_combout\);

-- Location: FF_X13_Y63_N13
\TheParToI2s|BclkCtr[2]~DUPLICATE\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \TheParToI2s|Selector7~1_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheParToI2s|BclkCtr[2]~DUPLICATE_q\);

-- Location: FF_X16_Y65_N20
\TheParToI2s|LastValidDL[1]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	asdata => \TheI2sToPar|D\(1),
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \TheI2sToPar|ValL~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheParToI2s|LastValidDL\(1));

-- Location: FF_X16_Y65_N59
\TheParToI2s|LastValidDL[3]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	asdata => \TheI2sToPar|D\(3),
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \TheI2sToPar|ValL~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheParToI2s|LastValidDL\(3));

-- Location: FF_X16_Y65_N5
\TheParToI2s|LastValidDL[9]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	asdata => \TheI2sToPar|D\(9),
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \TheI2sToPar|ValL~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheParToI2s|LastValidDL\(9));

-- Location: FF_X16_Y65_N56
\TheParToI2s|LastValidDL[11]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	asdata => \TheI2sToPar|D\(11),
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \TheI2sToPar|ValL~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheParToI2s|LastValidDL\(11));

-- Location: LABCELL_X16_Y65_N54
\TheParToI2s|Mux1~2\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheParToI2s|Mux1~2_combout\ = ( \TheParToI2s|LastValidDL\(11) & ( \TheParToI2s|BclkCtr[3]~DUPLICATE_q\ & ( (\TheParToI2s|BclkCtr\(1)) # (\TheParToI2s|LastValidDL\(9)) ) ) ) # ( !\TheParToI2s|LastValidDL\(11) & ( \TheParToI2s|BclkCtr[3]~DUPLICATE_q\ & ( 
-- (\TheParToI2s|LastValidDL\(9) & !\TheParToI2s|BclkCtr\(1)) ) ) ) # ( \TheParToI2s|LastValidDL\(11) & ( !\TheParToI2s|BclkCtr[3]~DUPLICATE_q\ & ( (!\TheParToI2s|BclkCtr\(1) & (\TheParToI2s|LastValidDL\(1))) # (\TheParToI2s|BclkCtr\(1) & 
-- ((\TheParToI2s|LastValidDL\(3)))) ) ) ) # ( !\TheParToI2s|LastValidDL\(11) & ( !\TheParToI2s|BclkCtr[3]~DUPLICATE_q\ & ( (!\TheParToI2s|BclkCtr\(1) & (\TheParToI2s|LastValidDL\(1))) # (\TheParToI2s|BclkCtr\(1) & ((\TheParToI2s|LastValidDL\(3)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101010100110011010101010011001100001111000000000000111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheParToI2s|ALT_INV_LastValidDL\(1),
	datab => \TheParToI2s|ALT_INV_LastValidDL\(3),
	datac => \TheParToI2s|ALT_INV_LastValidDL\(9),
	datad => \TheParToI2s|ALT_INV_BclkCtr\(1),
	datae => \TheParToI2s|ALT_INV_LastValidDL\(11),
	dataf => \TheParToI2s|ALT_INV_BclkCtr[3]~DUPLICATE_q\,
	combout => \TheParToI2s|Mux1~2_combout\);

-- Location: FF_X16_Y65_N47
\TheParToI2s|LastValidDL[13]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	asdata => \TheI2sToPar|D\(13),
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \TheI2sToPar|ValL~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheParToI2s|LastValidDL\(13));

-- Location: LABCELL_X16_Y65_N27
\TheParToI2s|LastValidDL[5]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheParToI2s|LastValidDL[5]~feeder_combout\ = ( \TheI2sToPar|D\(5) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \TheI2sToPar|ALT_INV_D\(5),
	combout => \TheParToI2s|LastValidDL[5]~feeder_combout\);

-- Location: FF_X16_Y65_N29
\TheParToI2s|LastValidDL[5]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \TheParToI2s|LastValidDL[5]~feeder_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	ena => \TheI2sToPar|ValL~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheParToI2s|LastValidDL\(5));

-- Location: FF_X16_Y65_N38
\TheParToI2s|LastValidDL[15]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	asdata => \TheI2sToPar|D\(15),
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \TheI2sToPar|ValL~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheParToI2s|LastValidDL\(15));

-- Location: FF_X16_Y65_N26
\TheParToI2s|LastValidDL[7]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	asdata => \TheI2sToPar|D\(7),
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \TheI2sToPar|ValL~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheParToI2s|LastValidDL\(7));

-- Location: LABCELL_X16_Y65_N36
\TheParToI2s|Mux1~3\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheParToI2s|Mux1~3_combout\ = ( \TheParToI2s|LastValidDL\(15) & ( \TheParToI2s|LastValidDL\(7) & ( ((!\TheParToI2s|BclkCtr[3]~DUPLICATE_q\ & ((\TheParToI2s|LastValidDL\(5)))) # (\TheParToI2s|BclkCtr[3]~DUPLICATE_q\ & (\TheParToI2s|LastValidDL\(13)))) # 
-- (\TheParToI2s|BclkCtr\(1)) ) ) ) # ( !\TheParToI2s|LastValidDL\(15) & ( \TheParToI2s|LastValidDL\(7) & ( (!\TheParToI2s|BclkCtr[3]~DUPLICATE_q\ & (((\TheParToI2s|BclkCtr\(1)) # (\TheParToI2s|LastValidDL\(5))))) # (\TheParToI2s|BclkCtr[3]~DUPLICATE_q\ & 
-- (\TheParToI2s|LastValidDL\(13) & ((!\TheParToI2s|BclkCtr\(1))))) ) ) ) # ( \TheParToI2s|LastValidDL\(15) & ( !\TheParToI2s|LastValidDL\(7) & ( (!\TheParToI2s|BclkCtr[3]~DUPLICATE_q\ & (((\TheParToI2s|LastValidDL\(5) & !\TheParToI2s|BclkCtr\(1))))) # 
-- (\TheParToI2s|BclkCtr[3]~DUPLICATE_q\ & (((\TheParToI2s|BclkCtr\(1))) # (\TheParToI2s|LastValidDL\(13)))) ) ) ) # ( !\TheParToI2s|LastValidDL\(15) & ( !\TheParToI2s|LastValidDL\(7) & ( (!\TheParToI2s|BclkCtr\(1) & ((!\TheParToI2s|BclkCtr[3]~DUPLICATE_q\ & 
-- ((\TheParToI2s|LastValidDL\(5)))) # (\TheParToI2s|BclkCtr[3]~DUPLICATE_q\ & (\TheParToI2s|LastValidDL\(13))))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0001101100000000000110110101010100011011101010100001101111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheParToI2s|ALT_INV_BclkCtr[3]~DUPLICATE_q\,
	datab => \TheParToI2s|ALT_INV_LastValidDL\(13),
	datac => \TheParToI2s|ALT_INV_LastValidDL\(5),
	datad => \TheParToI2s|ALT_INV_BclkCtr\(1),
	datae => \TheParToI2s|ALT_INV_LastValidDL\(15),
	dataf => \TheParToI2s|ALT_INV_LastValidDL\(7),
	combout => \TheParToI2s|Mux1~3_combout\);

-- Location: FF_X16_Y65_N40
\TheParToI2s|LastValidDL[2]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	asdata => \TheI2sToPar|D\(2),
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \TheI2sToPar|ValL~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheParToI2s|LastValidDL\(2));

-- Location: LABCELL_X16_Y65_N42
\TheParToI2s|LastValidDL[0]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheParToI2s|LastValidDL[0]~feeder_combout\ = ( \TheI2sToPar|D\(0) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \TheI2sToPar|ALT_INV_D\(0),
	combout => \TheParToI2s|LastValidDL[0]~feeder_combout\);

-- Location: FF_X16_Y65_N44
\TheParToI2s|LastValidDL[0]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \TheParToI2s|LastValidDL[0]~feeder_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	ena => \TheI2sToPar|ValL~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheParToI2s|LastValidDL\(0));

-- Location: LABCELL_X17_Y65_N51
\TheParToI2s|LastValidDL[8]~feeder\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheParToI2s|LastValidDL[8]~feeder_combout\ = ( \TheI2sToPar|D\(8) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000011111111111111111111111111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataf => \TheI2sToPar|ALT_INV_D\(8),
	combout => \TheParToI2s|LastValidDL[8]~feeder_combout\);

-- Location: FF_X17_Y65_N52
\TheParToI2s|LastValidDL[8]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	d => \TheParToI2s|LastValidDL[8]~feeder_combout\,
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	ena => \TheI2sToPar|ValL~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheParToI2s|LastValidDL\(8));

-- Location: FF_X16_Y65_N23
\TheParToI2s|LastValidDL[10]\ : dffeas
-- pragma translate_off
GENERIC MAP (
	is_wysiwyg => "true",
	power_up => "low")
-- pragma translate_on
PORT MAP (
	clk => \PLL_50MHz_48MHz|GeneratePLLForSyn:AlteraPLL50to48_rtl|alterapll50to48_inst|altera_pll_i|outclk_wire[0]~CLKENA0_outclk\,
	asdata => \TheI2sToPar|D\(10),
	clrn => \inResetAsync~inputCLKENA0_outclk\,
	sload => VCC,
	ena => \TheI2sToPar|ValL~q\,
	devclrn => ww_devclrn,
	devpor => ww_devpor,
	q => \TheParToI2s|LastValidDL\(10));

-- Location: LABCELL_X16_Y65_N21
\TheParToI2s|Mux1~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheParToI2s|Mux1~0_combout\ = ( \TheParToI2s|LastValidDL\(10) & ( \TheParToI2s|BclkCtr\(1) & ( (\TheParToI2s|BclkCtr[3]~DUPLICATE_q\) # (\TheParToI2s|LastValidDL\(2)) ) ) ) # ( !\TheParToI2s|LastValidDL\(10) & ( \TheParToI2s|BclkCtr\(1) & ( 
-- (\TheParToI2s|LastValidDL\(2) & !\TheParToI2s|BclkCtr[3]~DUPLICATE_q\) ) ) ) # ( \TheParToI2s|LastValidDL\(10) & ( !\TheParToI2s|BclkCtr\(1) & ( (!\TheParToI2s|BclkCtr[3]~DUPLICATE_q\ & (\TheParToI2s|LastValidDL\(0))) # 
-- (\TheParToI2s|BclkCtr[3]~DUPLICATE_q\ & ((\TheParToI2s|LastValidDL\(8)))) ) ) ) # ( !\TheParToI2s|LastValidDL\(10) & ( !\TheParToI2s|BclkCtr\(1) & ( (!\TheParToI2s|BclkCtr[3]~DUPLICATE_q\ & (\TheParToI2s|LastValidDL\(0))) # 
-- (\TheParToI2s|BclkCtr[3]~DUPLICATE_q\ & ((\TheParToI2s|LastValidDL\(8)))) ) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0011001100001111001100110000111101010101000000000101010111111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheParToI2s|ALT_INV_LastValidDL\(2),
	datab => \TheParToI2s|ALT_INV_LastValidDL\(0),
	datac => \TheParToI2s|ALT_INV_LastValidDL\(8),
	datad => \TheParToI2s|ALT_INV_BclkCtr[3]~DUPLICATE_q\,
	datae => \TheParToI2s|ALT_INV_LastValidDL\(10),
	dataf => \TheParToI2s|ALT_INV_BclkCtr\(1),
	combout => \TheParToI2s|Mux1~0_combout\);

-- Location: LABCELL_X16_Y65_N12
\TheParToI2s|Selector10~1\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheParToI2s|Selector10~1_combout\ = ( !\TheParToI2s|BclkCtr\(0) & ( ((\TheParToI2s|Selector10~0_combout\ & ((!\TheParToI2s|BclkCtr[2]~DUPLICATE_q\ & ((\TheParToI2s|Mux1~0_combout\))) # (\TheParToI2s|BclkCtr[2]~DUPLICATE_q\ & 
-- (\TheParToI2s|Mux1~1_combout\))))) ) ) # ( \TheParToI2s|BclkCtr\(0) & ( ((\TheParToI2s|Selector10~0_combout\ & ((!\TheParToI2s|BclkCtr[2]~DUPLICATE_q\ & (\TheParToI2s|Mux1~2_combout\)) # (\TheParToI2s|BclkCtr[2]~DUPLICATE_q\ & 
-- ((\TheParToI2s|Mux1~3_combout\)))))) ) )

-- pragma translate_off
GENERIC MAP (
	extended_lut => "on",
	lut_mask => "0000000000000000000000000000000000011101000111010000110000111111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheParToI2s|ALT_INV_Mux1~1_combout\,
	datab => \TheParToI2s|ALT_INV_BclkCtr[2]~DUPLICATE_q\,
	datac => \TheParToI2s|ALT_INV_Mux1~2_combout\,
	datad => \TheParToI2s|ALT_INV_Mux1~3_combout\,
	datae => \TheParToI2s|ALT_INV_BclkCtr\(0),
	dataf => \TheParToI2s|ALT_INV_Selector10~0_combout\,
	datag => \TheParToI2s|ALT_INV_Mux1~0_combout\,
	combout => \TheParToI2s|Selector10~1_combout\);

-- Location: LABCELL_X13_Y64_N39
\TheParToI2s|oLrc~0\ : cyclonev_lcell_comb
-- Equation(s):
-- \TheParToI2s|oLrc~0_combout\ = (\TheParToI2s|State.FirstBitEmptyL~q\) # (\TheParToI2s|State.SendingL~q\)

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0101111101011111010111110101111101011111010111110101111101011111",
	shared_arith => "off")
-- pragma translate_on
PORT MAP (
	dataa => \TheParToI2s|ALT_INV_State.SendingL~q\,
	datac => \TheParToI2s|ALT_INV_State.FirstBitEmptyL~q\,
	combout => \TheParToI2s|oLrc~0_combout\);

-- Location: IOIBUF_X16_Y0_N1
\iSwitch[1]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_iSwitch(1),
	o => \iSwitch[1]~input_o\);

-- Location: IOIBUF_X8_Y0_N35
\iSwitch[2]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_iSwitch(2),
	o => \iSwitch[2]~input_o\);

-- Location: IOIBUF_X4_Y0_N52
\iSwitch[3]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_iSwitch(3),
	o => \iSwitch[3]~input_o\);

-- Location: IOIBUF_X2_Y0_N41
\iSwitch[4]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_iSwitch(4),
	o => \iSwitch[4]~input_o\);

-- Location: IOIBUF_X16_Y0_N18
\iSwitch[5]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_iSwitch(5),
	o => \iSwitch[5]~input_o\);

-- Location: IOIBUF_X4_Y0_N35
\iSwitch[6]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_iSwitch(6),
	o => \iSwitch[6]~input_o\);

-- Location: IOIBUF_X4_Y0_N1
\iSwitch[7]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_iSwitch(7),
	o => \iSwitch[7]~input_o\);

-- Location: IOIBUF_X4_Y0_N18
\iSwitch[8]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_iSwitch(8),
	o => \iSwitch[8]~input_o\);

-- Location: IOIBUF_X2_Y0_N58
\iSwitch[9]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_iSwitch(9),
	o => \iSwitch[9]~input_o\);

-- Location: IOIBUF_X36_Y0_N18
\inButton[1]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_inButton(1),
	o => \inButton[1]~input_o\);

-- Location: IOIBUF_X40_Y0_N1
\inButton[2]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_inButton(2),
	o => \inButton[2]~input_o\);

-- Location: IOIBUF_X40_Y0_N18
\inButton[3]~input\ : cyclonev_io_ibuf
-- pragma translate_off
GENERIC MAP (
	bus_hold => "false",
	simulate_z_as => "z")
-- pragma translate_on
PORT MAP (
	i => ww_inButton(3),
	o => \inButton[3]~input_o\);

-- Location: LABCELL_X30_Y6_N3
\~QUARTUS_CREATED_GND~I\ : cyclonev_lcell_comb
-- Equation(s):

-- pragma translate_off
GENERIC MAP (
	extended_lut => "off",
	lut_mask => "0000000000000000000000000000000000000000000000000000000000000000",
	shared_arith => "off")
-- pragma translate_on
;


pll_reconfig_inst_tasks : altera_pll_reconfig_tasks
-- pragma translate_off
GENERIC MAP (
      number_of_fplls => 1);
-- pragma translate_on
END structure;


