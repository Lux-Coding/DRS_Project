--------------------------------------------------------------------------------
-- Title       : DDS sine wave generator
-- Project     : FPGA Based Digital Signal Processing
--               FH OÖ Hagenberg/HSD, SCD5
--------------------------------------------------------------------------------
-- RevCtrl     : $Id: DspDds-e.vhd 716 2017-11-12 16:57:46Z mroland $
-- Authors     : Markus Pfaff, Linz/Austria, Copyright (c) 2003-2005
--               Michael Roland, Hagenberg/Austria, Copyright (c) 2011-2017
--------------------------------------------------------------------------------
-- Description : 
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
-- Useful with some synthesis tools only. See architecture Rtl for more details.
-- use ieee.math_real.all;

-- fixed_pkg resides in the library ieee since VHDL-2008 (QuestaSim backports
-- this to VHDL-93 too). However, Quartus (as of version 13.0sp1) still does
-- not have native support for ieee.fixed_pkg. Therefore, we provide the
-- VHDL-93 compatibility versions as part of this excercise. These must be
-- compiled into the are located in the library ieee_proposed. Include them in
-- your Config.tcl and don't forget to set the ExtraLibraries and TargetLibrary
-- parameters to compile them into the right library (ieee_proposed) with fhlow.
library ieee_proposed;
use ieee_proposed.fixed_pkg.all;
use ieee_proposed.fixed_float_types.all;
-- In future (when both QuestaSim and Quartus support the VHDL-2008
-- ieee.fixed_pkg) simply use:
--use ieee.fixed_float_types.all;
--use ieee.fixed_pkg.all;

use work.Global.all;

entity DspDds is
  
  generic (
    gClkFrequency            : natural       := cDefaultClkFrequency;
    gAudioBitWidth           : natural       := cDefaultAudioBitWidth;

    -- How many bits does the phase register have?
    gPhaseResolution         : natural       := 20;

    -- How many bits of the phase register will be dithered?
    -- Should be gPhaseResolution-LogDualis(gWaveTable'length)
    -- Unfortunately this is not a globally static expression so we have
    -- express this via a literal.
    gNrOfPhaseDitherBits     : natural       := 8;

    -- How many bits do the waveform ROM table entries have?
    gWaveTableBitWidth       : natural       := 14;

    -- Precalculated waveform ROM table entries
    -- The values of the wave table are given for the first quadrant of
    -- the sine function. For more details see the paper from Martin
    -- Pechanec: "Output Spectrum of a Direct Digital Synthesizer".
    -- Can be found under the filename Dds.pdf on the internet.
   gWaveTable               : aSetOfFactors := (
	0.000766990318742704,
	0.0023009691514258,
	0.00383494256970623,
	0.00536890696399634,
	0.00690285872472976,
	0.0084367942423698,
	0.00997070990741803,
	0.0115046021104227,
	0.0130384672419873,
	0.0145723016927791,
	0.0161061018535373,
	0.0176398641150821,
	0.0191735848683226,
	0.0207072605042659,
	0.022240887414025,
	0.0237744619888276,
	0.0253079806200246,
	0.0268414396990985,
	0.0283748356176721,
	0.0299081647675166,
	0.0314414235405603,
	0.0329746083288973,
	0.0345077155247957,
	0.0360407415207062,
	0.0375736827092705,
	0.0391065354833299,
	0.0406392962359337,
	0.0421719613603479,
	0.0437045272500634,
	0.0452369902988046,
	0.0467693469005379,
	0.0483015934494801,
	0.0498337263401073,
	0.0513657419671626,
	0.0528976367256653,
	0.0544294070109191,
	0.0559610492185206,
	0.0574925597443676,
	0.0590239349846679,
	0.0605551713359478,
	0.0620862651950601,
	0.0636172129591931,
	0.0651480110258788,
	0.0666786557930016,
	0.0682091436588063,
	0.0697394710219073,
	0.0712696342812964,
	0.0727996298363517,
	0.0743294540868458,
	0.0758591034329544,
	0.077388574275265,
	0.0789178630147849,
	0.08044696605295,
	0.0819758797916331,
	0.0835046006331524,
	0.0850331249802803,
	0.0865614492362512,
	0.0880895698047705,
	0.089617483090023,
	0.091145185496681,
	0.0926726734299133,
	0.0941999432953932,
	0.0957269914993072,
	0.0972538144483633,
	0.0987804085497996,
	0.100306770211393,
	0.101832895841467,
	0.1033587818489,
	0.104884424643135,
	0.106409820634188,
	0.107934966232654,
	0.109459857849718,
	0.110984491897163,
	0.112508864787379,
	0.114032972933367,
	0.115556812748755,
	0.117080380647801,
	0.118603673045401,
	0.120126686357102,
	0.121649416999106,
	0.12317186138828,
	0.124694015942168,
	0.12621587707899,
	0.127737441217662,
	0.129258704777796,
	0.130779664179712,
	0.132300315844445,
	0.133820656193755,
	0.135340681650134,
	0.136860388636816,
	0.138379773577784,
	0.139898832897777,
	0.141417563022303,
	0.142935960377643,
	0.14445402139086,
	0.145971742489812,
	0.147489120103154,
	0.149006150660348,
	0.150522830591677,
	0.152039156328246,
	0.153555124301993,
	0.155070730945701,
	0.156585972692998,
	0.158100845978377,
	0.159615347237193,
	0.161129472905679,
	0.16264321942095,
	0.164156583221016,
	0.165669560744784,
	0.167182148432073,
	0.168694342723617,
	0.170206140061078,
	0.17171753688705,
	0.17322852964507,
	0.174739114779627,
	0.176249288736168,
	0.177759047961107,
	0.179268388901836,
	0.180777308006729,
	0.182285801725153,
	0.183793866507478,
	0.185301498805082,
	0.186808695070359,
	0.188315451756732,
	0.189821765318656,
	0.191327632211631,
	0.192833048892205,
	0.194338011817989,
	0.195842517447658,
	0.197346562240966,
	0.19885014265875,
	0.20035325516294,
	0.201855896216568,
	0.203358062283773,
	0.204859749829814,
	0.206360955321076,
	0.207861675225075,
	0.209361906010474,
	0.210861644147085,
	0.212360886105878,
	0.213859628358994,
	0.215357867379746,
	0.216855599642633,
	0.218352821623346,
	0.219849529798779,
	0.221345720647031,
	0.222841390647421,
	0.224336536280494,
	0.225831154028026,
	0.227325240373039,
	0.228818791799802,
	0.230311804793845,
	0.231804275841965,
	0.233296201432232,
	0.234787578054001,
	0.23627840219792,
	0.237768670355934,
	0.2392583790213,
	0.240747524688588,
	0.242236103853696,
	0.243724113013852,
	0.245211548667628,
	0.246698407314942,
	0.248184685457075,
	0.249670379596669,
	0.251155486237742,
	0.252640001885696,
	0.254123923047321,
	0.255607246230807,
	0.257089967945753,
	0.25857208470317,
	0.260053593015495,
	0.261534489396596,
	0.263014770361779,
	0.264494432427802,
	0.265973472112876,
	0.267451885936678,
	0.268929670420357,
	0.270406822086545,
	0.27188333745936,
	0.273359213064419,
	0.274834445428844,
	0.276309031081271,
	0.277782966551858,
	0.279256248372291,
	0.280728873075797,
	0.282200837197148,
	0.283672137272668,
	0.285142769840249,
	0.286612731439348,
	0.288082018611004,
	0.289550627897843,
	0.291018555844085,
	0.292485798995554,
	0.293952353899685,
	0.295418217105532,
	0.296883385163778,
	0.298347854626741,
	0.299811622048383,
	0.301274683984318,
	0.302737036991819,
	0.304198677629829,
	0.305659602458966,
	0.307119808041533,
	0.308579290941525,
	0.310038047724638,
	0.311496074958276,
	0.31295336921156,
	0.314409927055337,
	0.315865745062184,
	0.317320819806422,
	0.318775147864119,
	0.3202287258131,
	0.321681550232957,
	0.323133617705052,
	0.324584924812532,
	0.32603546814033,
	0.327485244275178,
	0.328934249805612,
	0.330382481321983,
	0.331829935416461,
	0.333276608683048,
	0.334722497717581,
	0.336167599117745,
	0.337611909483075,
	0.33905542541497,
	0.340498143516697,
	0.341940060393402,
	0.343381172652115,
	0.344821476901759,
	0.34626096975316,
	0.347699647819051,
	0.349137507714085,
	0.350574546054838,
	0.352010759459819,
	0.353446144549481,
	0.354880697946223,
	0.356314416274402,
	0.357747296160342,
	0.359179334232337,
	0.360610527120662,
	0.362040871457584,
	0.363470363877364,
	0.364899001016267,
	0.366326779512574,
	0.367753696006582,
	0.36917974714062,
	0.370604929559052,
	0.372029239908285,
	0.37345267483678,
	0.374875230995058,
	0.376296905035705,
	0.377717693613386,
	0.379137593384847,
	0.380556601008929,
	0.381974713146567,
	0.383391926460809,
	0.384808237616813,
	0.386223643281863,
	0.387638140125373,
	0.389051724818894,
	0.390464394036127,
	0.391876144452922,
	0.393286972747296,
	0.394696875599434,
	0.396105849691696,
	0.397513891708632,
	0.398920998336983,
	0.40032716626569,
	0.401732392185905,
	0.403136672790995,
	0.404540004776553,
	0.405942384840403,
	0.407343809682608,
	0.408744276005481,
	0.41014378051359,
	0.411542319913765,
	0.412939890915108,
	0.414336490228999,
	0.415732114569105,
	0.417126760651388,
	0.41852042519411,
	0.419913104917844,
	0.42130479654548,
	0.422695496802233,
	0.424085202415652,
	0.425473910115624,
	0.426861616634386,
	0.428248318706532,
	0.429634013069016,
	0.431018696461167,
	0.43240236562469,
	0.433785017303679,
	0.435166648244619,
	0.436547255196401,
	0.437926834910323,
	0.4393053841401,
	0.440682899641873,
	0.442059378174215,
	0.443434816498138,
	0.444809211377105,
	0.44618255957703,
	0.447554857866293,
	0.448926103015743,
	0.450296291798709,
	0.451665420991003,
	0.453033487370932,
	0.454400487719304,
	0.455766418819435,
	0.457131277457157,
	0.458495060420826,
	0.45985776450133,
	0.461219386492092,
	0.462579923189087,
	0.463939371390839,
	0.465297727898435,
	0.466654989515531,
	0.46801115304836,
	0.469366215305738,
	0.470720173099072,
	0.472073023242369,
	0.473424762552242,
	0.474775387847917,
	0.476124895951244,
	0.477473283686698,
	0.478820547881394,
	0.480166685365088,
	0.48151169297019,
	0.482855567531766,
	0.484198305887549,
	0.485539904877947,
	0.486880361346047,
	0.488219672137627,
	0.489557834101157,
	0.490894844087815,
	0.492230698951486,
	0.493565395548775,
	0.494898930739011,
	0.496231301384258,
	0.497562504349319,
	0.498892536501745,
	0.500221394711841,
	0.501549075852675,
	0.502875576800087,
	0.50420089443269,
	0.505525025631885,
	0.506847967281863,
	0.508169716269615,
	0.509490269484936,
	0.510809623820439,
	0.512127776171555,
	0.513444723436543,
	0.514760462516501,
	0.516074990315367,
	0.517388303739929,
	0.518700399699835,
	0.520011275107596,
	0.521320926878596,
	0.522629351931097,
	0.523936547186248,
	0.525242509568095,
	0.526547236003579,
	0.527850723422555,
	0.529152968757791,
	0.530453968944976,
	0.531753720922733,
	0.533052221632619,
	0.534349468019138,
	0.535645457029741,
	0.536940185614843,
	0.538233650727822,
	0.539525849325029,
	0.540816778365797,
	0.542106434812444,
	0.543394815630285,
	0.544681917787635,
	0.545967738255818,
	0.547252274009174,
	0.548535522025067,
	0.549817479283891,
	0.551098142769075,
	0.552377509467096,
	0.553655576367479,
	0.55493234046281,
	0.55620779874874,
	0.557481948223992,
	0.558754785890368,
	0.56002630875276,
	0.561296513819151,
	0.562565398100626,
	0.563832958611378,
	0.565099192368714,
	0.566364096393064,
	0.567627667707986,
	0.568889903340176,
	0.57015080031947,
	0.571410355678857,
	0.572668566454481,
	0.573925429685651,
	0.575180942414845,
	0.576435101687722,
	0.577687904553123,
	0.578939348063082,
	0.580189429272832,
	0.58143814524081,
	0.582685493028668,
	0.583931469701276,
	0.58517607232673,
	0.58641929797636,
	0.587661143724737,
	0.588901606649676,
	0.590140683832249,
	0.591378372356787,
	0.592614669310891,
	0.593849571785434,
	0.59508307687457,
	0.596315181675744,
	0.597545883289693,
	0.598775178820459,
	0.600003065375389,
	0.601229540065149,
	0.602454600003724,
	0.60367824230843,
	0.60490046409992,
	0.606121262502186,
	0.607340634642573,
	0.608558577651779,
	0.609775088663868,
	0.610990164816272,
	0.612203803249798,
	0.613416001108639,
	0.614626755540375,
	0.615836063695985,
	0.61704392272985,
	0.61825032979976,
	0.619455282066924,
	0.620658776695972,
	0.621860810854965,
	0.623061381715401,
	0.624260486452221,
	0.625458122243814,
	0.626654286272029,
	0.627848975722177,
	0.629042187783036,
	0.630233919646864,
	0.631424168509402,
	0.632612931569877,
	0.633800206031017,
	0.634985989099049,
	0.636170277983712,
	0.637353069898259,
	0.638534362059467,
	0.63971415168764,
	0.640892436006621,
	0.642069212243792,
	0.643244477630086,
	0.644418229399988,
	0.645590464791549,
	0.646761181046384,
	0.647930375409685,
	0.649098045130226,
	0.650264187460366,
	0.65142879965606,
	0.652591878976862,
	0.653753422685936,
	0.654913428050056,
	0.656071892339618,
	0.657228812828643,
	0.658384186794785,
	0.659538011519339,
	0.660690284287242,
	0.661841002387087,
	0.662990163111121,
	0.66413776375526,
	0.665283801619087,
	0.666428274005865,
	0.66757117822254,
	0.668712511579748,
	0.669852271391821,
	0.670990454976794,
	0.672127059656412,
	0.673262082756133,
	0.674395521605139,
	0.675527373536339,
	0.676657635886375,
	0.677786305995631,
	0.678913381208238,
	0.680038858872079,
	0.681162736338795,
	0.682285010963795,
	0.683405680106259,
	0.684524741129142,
	0.685642191399187,
	0.686758028286926,
	0.687872249166686,
	0.688984851416597,
	0.6900958324186,
	0.691205189558448,
	0.692312920225718,
	0.693419021813812,
	0.694523491719965,
	0.695626327345255,
	0.696727526094601,
	0.697827085376777,
	0.698925002604414,
	0.700021275194006,
	0.701115900565919,
	0.702208876144392,
	0.703300199357549,
	0.7043898676374,
	0.705477878419852,
	0.70656422914471,
	0.707648917255684,
	0.708731940200401,
	0.709813295430401,
	0.710892980401152,
	0.71197099257205,
	0.713047329406429,
	0.714121988371565,
	0.71519496693868,
	0.716266262582953,
	0.717335872783522,
	0.71840379502349,
	0.719470026789933,
	0.720534565573905,
	0.721597408870444,
	0.722658554178576,
	0.723717999001323,
	0.724775740845711,
	0.72583177722277,
	0.726886105647545,
	0.727938723639099,
	0.728989628720519,
	0.730038818418926,
	0.731086290265474,
	0.732132041795361,
	0.733176070547833,
	0.734218374066188,
	0.735258949897787,
	0.736297795594053,
	0.737334908710483,
	0.738370286806649,
	0.739403927446206,
	0.740435828196898,
	0.741465986630563,
	0.742494400323139,
	0.743521066854669,
	0.744545983809307,
	0.745569148775325,
	0.746590559345117,
	0.747610213115205,
	0.748628107686245,
	0.749644240663033,
	0.750658609654511,
	0.751671212273768,
	0.752682046138055,
	0.753691108868781,
	0.754698398091525,
	0.755703911436036,
	0.756707646536246,
	0.757709601030268,
	0.758709772560407,
	0.759708158773163,
	0.760704757319237,
	0.761699565853535,
	0.762692582035178,
	0.763683803527502,
	0.764673227998067,
	0.765660853118662,
	0.76664667656531,
	0.767630696018273,
	0.768612909162058,
	0.769593313685423,
	0.770571907281381,
	0.771548687647206,
	0.772523652484441,
	0.773496799498899,
	0.774468126400671,
	0.775437630904131,
	0.77640531072794,
	0.777371163595056,
	0.778335187232733,
	0.77929737937253,
	0.780257737750317,
	0.781216260106276,
	0.782172944184913,
	0.783127787735057,
	0.78408078850987,
	0.785031944266848,
	0.78598125276783,
	0.786928711779002,
	0.7878743190709,
	0.78881807241842,
	0.789759969600819,
	0.790700008401722,
	0.791638186609126,
	0.792574502015408,
	0.793508952417327,
	0.794441535616031,
	0.795372249417061,
	0.796301091630359,
	0.797228060070269,
	0.798153152555544,
	0.799076366909352,
	0.799997700959282,
	0.800917152537344,
	0.801834719479981,
	0.802750399628069,
	0.803664190826924,
	0.804576090926307,
	0.805486097780429,
	0.806394209247956,
	0.807300423192014,
	0.808204737480195,
	0.809107149984558,
	0.810007658581641,
	0.81090626115246,
	0.811802955582515,
	0.812697739761799,
	0.813590611584799,
	0.814481568950499,
	0.815370609762391,
	0.816257731928477,
	0.817142933361273,
	0.818026211977813,
	0.818907565699659,
	0.819786992452899,
	0.820664490168157,
	0.821540056780597,
	0.822413690229926,
	0.8232853884604,
	0.824155149420829,
	0.82502297106458,
	0.825888851349587,
	0.826752788238349,
	0.827614779697938,
	0.828474823700007,
	0.829332918220788,
	0.830189061241102,
	0.831043250746362,
	0.831895484726578,
	0.832745761176359,
	0.833594078094925,
	0.834440433486103,
	0.835284825358337,
	0.836127251724692,
	0.836967710602857,
	0.837806200015151,
	0.838642717988527,
	0.839477262554579,
	0.840309831749541,
	0.841140423614298,
	0.841969036194388,
	0.842795667540004,
	0.843620315706004,
	0.844442978751911,
	0.845263654741918,
	0.846082341744897,
	0.846899037834397,
	0.847713741088654,
	0.848526449590593,
	0.849337161427831,
	0.850145874692685,
	0.850952587482176,
	0.851757297898029,
	0.852560004046684,
	0.853360704039295,
	0.854159395991739,
	0.854956078024615,
	0.855750748263254,
	0.85654340483772,
	0.857334045882816,
	0.858122669538086,
	0.858909273947824,
	0.859693857261073,
	0.860476417631632,
	0.861256953218062,
	0.862035462183687,
	0.8628119426966,
	0.863586392929668,
	0.864358811060534,
	0.865129195271624,
	0.865897543750149,
	0.866663854688111,
	0.867428126282307,
	0.868190356734331,
	0.868950544250582,
	0.869708687042266,
	0.870464783325398,
	0.871218831320811,
	0.871970829254158,
	0.872720775355914,
	0.873468667861385,
	0.874214505010706,
	0.874958285048852,
	0.875700006225635,
	0.876439666795714,
	0.877177265018596,
	0.877912799158642,
	0.878646267485068,
	0.879377668271953,
	0.88010699979824,
	0.880834260347742,
	0.881559448209144,
	0.882282561676009,
	0.883003599046781,
	0.88372255862479,
	0.884439438718254,
	0.885154237640285,
	0.885866953708893,
	0.886577585246987,
	0.887286130582383,
	0.887992588047806,
	0.888696955980892,
	0.889399232724196,
	0.890099416625192,
	0.890797506036282,
	0.891493499314791,
	0.892187394822982,
	0.892879190928052,
	0.893568886002136,
	0.894256478422316,
	0.894941966570621,
	0.89562534883403,
	0.89630662360448,
	0.896985789278864,
	0.897662844259041,
	0.898337786951834,
	0.899010615769039,
	0.899681329127424,
	0.900349925448736,
	0.901016403159702,
	0.901680760692038,
	0.902342996482444,
	0.903003108972617,
	0.903661096609248,
	0.904316957844028,
	0.904970691133653,
	0.905622294939825,
	0.906271767729258,
	0.906919107973678,
	0.907564314149833,
	0.908207384739489,
	0.908848318229439,
	0.909487113111505,
	0.910123767882542,
	0.910758281044438,
	0.911390651104122,
	0.912020876573568,
	0.912648955969794,
	0.913274887814868,
	0.913898670635912,
	0.914520302965105,
	0.915139783339685,
	0.915757110301957,
	0.916372282399289,
	0.916985298184123,
	0.917596156213973,
	0.918204855051431,
	0.91881139326417,
	0.919415769424947,
	0.920017982111607,
	0.920618029907084,
	0.921215911399409,
	0.921811625181708,
	0.92240516985221,
	0.922996544014246,
	0.923585746276257,
	0.924172775251791,
	0.924757629559514,
	0.925340307823206,
	0.92592080867177,
	0.926499130739231,
	0.92707527266474,
	0.927649233092581,
	0.928221010672169,
	0.928790604058057,
	0.929358011909935,
	0.92992323289264,
	0.93048626567615,
	0.931047108935595,
	0.931605761351258,
	0.932162221608574,
	0.93271648839814,
	0.933268560415712,
	0.933818436362211,
	0.934366114943726,
	0.934911594871516,
	0.935454874862015,
	0.935995953636831,
	0.936534829922755,
	0.937071502451759,
	0.937605969961,
	0.938138231192824,
	0.93866828489477,
	0.93919612981957,
	0.939721764725153,
	0.940245188374651,
	0.940766399536396,
	0.941285396983929,
	0.941802179495998,
	0.942316745856564,
	0.942829094854803,
	0.943339225285108,
	0.943847135947093,
	0.944352825645595,
	0.944856293190677,
	0.945357537397632,
	0.945856557086984,
	0.946353351084491,
	0.946847918221148,
	0.947340257333192,
	0.947830367262101,
	0.948318246854599,
	0.948803894962658,
	0.949287310443502,
	0.949768492159607,
	0.950247438978705,
	0.95072414977379,
	0.951198623423113,
	0.951670858810194,
	0.952140854823816,
	0.952608610358033,
	0.953074124312172,
	0.953537395590833,
	0.953998423103895,
	0.954457205766514,
	0.954913742499131,
	0.95536803222747,
	0.955820073882545,
	0.956269866400658,
	0.956717408723403,
	0.95716269979767,
	0.957605738575646,
	0.958046524014819,
	0.958485055077976,
	0.958921330733213,
	0.959355349953931,
	0.95978711171884,
	0.960216615011963,
	0.960643858822639,
	0.961068842145519,
	0.961491563980579,
	0.961912023333112,
	0.962330219213737,
	0.962746150638399,
	0.963159816628371,
	0.963571216210257,
	0.963980348415994,
	0.964387212282854,
	0.964791806853448,
	0.965194131175725,
	0.965594184302977,
	0.965991965293841,
	0.966387473212299,
	0.966780707127683,
	0.967171666114677,
	0.967560349253314,
	0.967946755628988,
	0.968330884332445,
	0.968712734459795,
	0.969092305112506,
	0.969469595397413,
	0.969844604426715,
	0.970217331317979,
	0.970587775194144,
	0.970955935183518,
	0.971321810419786,
	0.971685400042009,
	0.972046703194623,
	0.97240571902745,
	0.972762446695689,
	0.973116885359925,
	0.973469034186131,
	0.973818892345666,
	0.97416645901528,
	0.974511733377116,
	0.974854714618708,
	0.97519540193299,
	0.975533794518291,
	0.975869891578341,
	0.976203692322271,
	0.976535195964614,
	0.976864401725313,
	0.977191308829712,
	0.977515916508569,
	0.97783822399805,
	0.978158230539735,
	0.978475935380617,
	0.978791337773106,
	0.979104436975029,
	0.979415232249635,
	0.979723722865591,
	0.98002990809699,
	0.980333787223348,
	0.980635359529608,
	0.980934624306142,
	0.98123158084875,
	0.981526228458665,
	0.981818566442552,
	0.982108594112514,
	0.982396310786085,
	0.982681715786241,
	0.982964808441396,
	0.983245588085407,
	0.983524054057571,
	0.983800205702632,
	0.984074042370776,
	0.984345563417642,
	0.984614768204313,
	0.984881656097324,
	0.985146226468662,
	0.985408478695768,
	0.985668412161538,
	0.985926026254321,
	0.986181320367928,
	0.986434293901627,
	0.986684946260147,
	0.986933276853678,
	0.987179285097874,
	0.987422970413855,
	0.987664332228206,
	0.987903369972978,
	0.988140083085693,
	0.988374471009341,
	0.988606533192386,
	0.988836269088764,
	0.989063678157882,
	0.989288759864625,
	0.989511513679355,
	0.989731939077911,
	0.989950035541609,
	0.990165802557248,
	0.990379239617108,
	0.99059034621895,
	0.99079912186602,
	0.991005566067049,
	0.991209678336254,
	0.991411458193339,
	0.991610905163495,
	0.991808018777406,
	0.992002798571245,
	0.992195244086674,
	0.992385354870852,
	0.992573130476429,
	0.992758570461551,
	0.99294167438986,
	0.993122441830496,
	0.993300872358093,
	0.993476965552789,
	0.993650721000219,
	0.99382213829152,
	0.993991217023329,
	0.99415795679779,
	0.994322357222546,
	0.994484417910748,
	0.994644138481051,
	0.994801518557617,
	0.994956557770116,
	0.995109255753726,
	0.995259612149133,
	0.995407626602535,
	0.995553298765638,
	0.995696628295664,
	0.995837614855342,
	0.995976258112918,
	0.996112557742151,
	0.996246513422316,
	0.9963781248382,
	0.996507391680111,
	0.99663431364387,
	0.996758890430818,
	0.996881121747814,
	0.997001007307235,
	0.99711854682698,
	0.997233740030466,
	0.997346586646633,
	0.997457086409942,
	0.997565239060376,
	0.997671044343441,
	0.997774502010168,
	0.99787561181711,
	0.997974373526347,
	0.998070786905482,
	0.998164851727646,
	0.998256567771495,
	0.998345934821212,
	0.998432952666508,
	0.998517621102622,
	0.99859993993032,
	0.998679908955899,
	0.998757527991183,
	0.998832796853528,
	0.998905715365818,
	0.99897628335647,
	0.999044500659429,
	0.999110367114175,
	0.999173882565716,
	0.999235046864596,
	0.999293859866888,
	0.999350321434199,
	0.999404431433671,
	0.999456189737977,
	0.999505596225325,
	0.999552650779457,
	0.999597353289648,
	0.99963970365071,
	0.999679701762988,
	0.999717347532362,
	0.999752640870249,
	0.999785581693599,
	0.9998161699249,
	0.999844405492175,
	0.999870288328983,
	0.999893818374418,
	0.999914995573113,
	0.999933819875236,
	0.99995029123649,
	0.999964409618118,
	0.999976174986898,
	0.999985587315143,
	0.999992646580707,
	0.999997352766978,
	0.999999705862882,
	0.999999705862882,
	0.999997352766978,
	0.999992646580707,
	0.999985587315143,
	0.999976174986898,
	0.999964409618118,
	0.99995029123649,
	0.999933819875236,
	0.999914995573113,
	0.999893818374418,
	0.999870288328983,
	0.999844405492175,
	0.9998161699249,
	0.999785581693599,
	0.999752640870249,
	0.999717347532362,
	0.999679701762988,
	0.99963970365071,
	0.999597353289648,
	0.999552650779457,
	0.999505596225325,
	0.999456189737977,
	0.999404431433671,
	0.999350321434199,
	0.999293859866888,
	0.999235046864596,
	0.999173882565716,
	0.999110367114175,
	0.999044500659429,
	0.99897628335647,
	0.998905715365818,
	0.998832796853528,
	0.998757527991183,
	0.998679908955899,
	0.99859993993032,
	0.998517621102622,
	0.998432952666508,
	0.998345934821212,
	0.998256567771495,
	0.998164851727646,
	0.998070786905482,
	0.997974373526347,
	0.99787561181711,
	0.997774502010168,
	0.997671044343441,
	0.997565239060376,
	0.997457086409942,
	0.997346586646633,
	0.997233740030466,
	0.99711854682698,
	0.997001007307235,
	0.996881121747814,
	0.996758890430818,
	0.99663431364387,
	0.996507391680111,
	0.9963781248382,
	0.996246513422316,
	0.996112557742151,
	0.995976258112918,
	0.995837614855342,
	0.995696628295664,
	0.995553298765638,
	0.995407626602535,
	0.995259612149133,
	0.995109255753726,
	0.994956557770116,
	0.994801518557617,
	0.994644138481051,
	0.994484417910748,
	0.994322357222546,
	0.99415795679779,
	0.993991217023329,
	0.99382213829152,
	0.993650721000219,
	0.993476965552789,
	0.993300872358093,
	0.993122441830496,
	0.99294167438986,
	0.992758570461551,
	0.992573130476429,
	0.992385354870852,
	0.992195244086674,
	0.992002798571245,
	0.991808018777406,
	0.991610905163495,
	0.991411458193339,
	0.991209678336254,
	0.991005566067049,
	0.99079912186602,
	0.99059034621895,
	0.990379239617108,
	0.990165802557248,
	0.989950035541609,
	0.989731939077911,
	0.989511513679355,
	0.989288759864625,
	0.989063678157882,
	0.988836269088764,
	0.988606533192386,
	0.988374471009341,
	0.988140083085693,
	0.987903369972978,
	0.987664332228206,
	0.987422970413855,
	0.987179285097874,
	0.986933276853678,
	0.986684946260147,
	0.986434293901627,
	0.986181320367928,
	0.985926026254321,
	0.985668412161538,
	0.985408478695768,
	0.985146226468662,
	0.984881656097324,
	0.984614768204313,
	0.984345563417642,
	0.984074042370776,
	0.983800205702632,
	0.983524054057571,
	0.983245588085407,
	0.982964808441396,
	0.982681715786241,
	0.982396310786085,
	0.982108594112513,
	0.981818566442552,
	0.981526228458665,
	0.98123158084875,
	0.980934624306142,
	0.980635359529608,
	0.980333787223348,
	0.98002990809699,
	0.979723722865591,
	0.979415232249635,
	0.979104436975029,
	0.978791337773106,
	0.978475935380617,
	0.978158230539735,
	0.97783822399805,
	0.977515916508569,
	0.977191308829712,
	0.976864401725313,
	0.976535195964614,
	0.976203692322271,
	0.975869891578341,
	0.975533794518291,
	0.97519540193299,
	0.974854714618708,
	0.974511733377116,
	0.97416645901528,
	0.973818892345666,
	0.973469034186131,
	0.973116885359925,
	0.972762446695689,
	0.97240571902745,
	0.972046703194623,
	0.971685400042009,
	0.971321810419786,
	0.970955935183518,
	0.970587775194144,
	0.970217331317979,
	0.969844604426715,
	0.969469595397413,
	0.969092305112506,
	0.968712734459795,
	0.968330884332445,
	0.967946755628988,
	0.967560349253314,
	0.967171666114677,
	0.966780707127683,
	0.966387473212299,
	0.965991965293841,
	0.965594184302977,
	0.965194131175725,
	0.964791806853448,
	0.964387212282854,
	0.963980348415994,
	0.963571216210257,
	0.963159816628371,
	0.962746150638399,
	0.962330219213737,
	0.961912023333112,
	0.961491563980579,
	0.961068842145519,
	0.960643858822639,
	0.960216615011963,
	0.95978711171884,
	0.959355349953931,
	0.958921330733213,
	0.958485055077976,
	0.958046524014818,
	0.957605738575646,
	0.95716269979767,
	0.956717408723403,
	0.956269866400658,
	0.955820073882545,
	0.95536803222747,
	0.95491374249913,
	0.954457205766513,
	0.953998423103894,
	0.953537395590833,
	0.953074124312172,
	0.952608610358033,
	0.952140854823816,
	0.951670858810194,
	0.951198623423113,
	0.95072414977379,
	0.950247438978705,
	0.949768492159607,
	0.949287310443502,
	0.948803894962658,
	0.948318246854599,
	0.947830367262101,
	0.947340257333192,
	0.946847918221148,
	0.946353351084491,
	0.945856557086984,
	0.945357537397632,
	0.944856293190677,
	0.944352825645595,
	0.943847135947093,
	0.943339225285108,
	0.942829094854803,
	0.942316745856564,
	0.941802179495998,
	0.941285396983929,
	0.940766399536396,
	0.940245188374651,
	0.939721764725153,
	0.93919612981957,
	0.93866828489477,
	0.938138231192824,
	0.937605969961,
	0.937071502451759,
	0.936534829922755,
	0.935995953636831,
	0.935454874862015,
	0.934911594871516,
	0.934366114943726,
	0.933818436362211,
	0.933268560415712,
	0.93271648839814,
	0.932162221608574,
	0.931605761351258,
	0.931047108935595,
	0.93048626567615,
	0.92992323289264,
	0.929358011909936,
	0.928790604058057,
	0.928221010672169,
	0.927649233092581,
	0.92707527266474,
	0.926499130739231,
	0.92592080867177,
	0.925340307823206,
	0.924757629559514,
	0.924172775251791,
	0.923585746276257,
	0.922996544014246,
	0.92240516985221,
	0.921811625181708,
	0.921215911399409,
	0.920618029907084,
	0.920017982111606,
	0.919415769424947,
	0.91881139326417,
	0.918204855051431,
	0.917596156213973,
	0.916985298184123,
	0.916372282399289,
	0.915757110301957,
	0.915139783339685,
	0.914520302965104,
	0.913898670635912,
	0.913274887814868,
	0.912648955969794,
	0.912020876573568,
	0.911390651104122,
	0.910758281044438,
	0.910123767882542,
	0.909487113111505,
	0.908848318229439,
	0.908207384739489,
	0.907564314149833,
	0.906919107973678,
	0.906271767729258,
	0.905622294939825,
	0.904970691133653,
	0.904316957844028,
	0.903661096609248,
	0.903003108972617,
	0.902342996482444,
	0.901680760692038,
	0.901016403159702,
	0.900349925448736,
	0.899681329127424,
	0.899010615769039,
	0.898337786951834,
	0.897662844259041,
	0.896985789278864,
	0.89630662360448,
	0.89562534883403,
	0.894941966570621,
	0.894256478422316,
	0.893568886002136,
	0.892879190928052,
	0.892187394822983,
	0.891493499314791,
	0.890797506036282,
	0.890099416625192,
	0.889399232724196,
	0.888696955980892,
	0.887992588047806,
	0.887286130582383,
	0.886577585246987,
	0.885866953708893,
	0.885154237640285,
	0.884439438718254,
	0.88372255862479,
	0.883003599046781,
	0.882282561676009,
	0.881559448209144,
	0.880834260347742,
	0.88010699979824,
	0.879377668271953,
	0.878646267485068,
	0.877912799158642,
	0.877177265018596,
	0.876439666795714,
	0.875700006225635,
	0.874958285048852,
	0.874214505010706,
	0.873468667861385,
	0.872720775355914,
	0.871970829254158,
	0.871218831320811,
	0.870464783325398,
	0.869708687042266,
	0.868950544250582,
	0.868190356734331,
	0.867428126282307,
	0.866663854688111,
	0.865897543750149,
	0.865129195271624,
	0.864358811060534,
	0.863586392929668,
	0.8628119426966,
	0.862035462183687,
	0.861256953218062,
	0.860476417631632,
	0.859693857261073,
	0.858909273947824,
	0.858122669538086,
	0.857334045882816,
	0.85654340483772,
	0.855750748263254,
	0.854956078024615,
	0.854159395991739,
	0.853360704039296,
	0.852560004046684,
	0.851757297898029,
	0.850952587482176,
	0.850145874692685,
	0.849337161427831,
	0.848526449590593,
	0.847713741088654,
	0.846899037834397,
	0.846082341744897,
	0.845263654741918,
	0.844442978751911,
	0.843620315706004,
	0.842795667540004,
	0.841969036194388,
	0.841140423614298,
	0.840309831749541,
	0.839477262554579,
	0.838642717988527,
	0.837806200015151,
	0.836967710602857,
	0.836127251724692,
	0.835284825358337,
	0.834440433486103,
	0.833594078094925,
	0.832745761176359,
	0.831895484726578,
	0.831043250746362,
	0.830189061241102,
	0.829332918220788,
	0.828474823700007,
	0.827614779697938,
	0.826752788238349,
	0.825888851349587,
	0.82502297106458,
	0.824155149420828,
	0.8232853884604,
	0.822413690229926,
	0.821540056780597,
	0.820664490168157,
	0.819786992452899,
	0.818907565699659,
	0.818026211977813,
	0.817142933361273,
	0.816257731928478,
	0.815370609762391,
	0.814481568950499,
	0.813590611584799,
	0.812697739761799,
	0.811802955582515,
	0.81090626115246,
	0.810007658581641,
	0.809107149984558,
	0.808204737480195,
	0.807300423192014,
	0.806394209247956,
	0.805486097780429,
	0.804576090926307,
	0.803664190826924,
	0.802750399628069,
	0.801834719479981,
	0.800917152537344,
	0.799997700959282,
	0.799076366909352,
	0.798153152555544,
	0.797228060070269,
	0.796301091630359,
	0.795372249417061,
	0.79444153561603,
	0.793508952417327,
	0.792574502015408,
	0.791638186609126,
	0.790700008401722,
	0.789759969600819,
	0.78881807241842,
	0.7878743190709,
	0.786928711779002,
	0.78598125276783,
	0.785031944266848,
	0.78408078850987,
	0.783127787735057,
	0.782172944184913,
	0.781216260106276,
	0.780257737750317,
	0.77929737937253,
	0.778335187232733,
	0.777371163595056,
	0.77640531072794,
	0.775437630904131,
	0.774468126400671,
	0.773496799498899,
	0.772523652484441,
	0.771548687647206,
	0.770571907281381,
	0.769593313685423,
	0.768612909162058,
	0.767630696018273,
	0.76664667656531,
	0.765660853118662,
	0.764673227998067,
	0.763683803527502,
	0.762692582035178,
	0.761699565853535,
	0.760704757319237,
	0.759708158773163,
	0.758709772560408,
	0.757709601030268,
	0.756707646536246,
	0.755703911436036,
	0.754698398091524,
	0.753691108868781,
	0.752682046138055,
	0.751671212273768,
	0.750658609654511,
	0.749644240663033,
	0.748628107686245,
	0.747610213115205,
	0.746590559345117,
	0.745569148775326,
	0.744545983809307,
	0.743521066854669,
	0.742494400323139,
	0.741465986630563,
	0.740435828196898,
	0.739403927446206,
	0.738370286806649,
	0.737334908710483,
	0.736297795594053,
	0.735258949897787,
	0.734218374066188,
	0.733176070547833,
	0.732132041795361,
	0.731086290265474,
	0.730038818418926,
	0.728989628720519,
	0.727938723639099,
	0.726886105647545,
	0.72583177722277,
	0.724775740845711,
	0.723717999001323,
	0.722658554178576,
	0.721597408870444,
	0.720534565573905,
	0.719470026789933,
	0.71840379502349,
	0.717335872783522,
	0.716266262582953,
	0.71519496693868,
	0.714121988371565,
	0.713047329406429,
	0.71197099257205,
	0.710892980401152,
	0.709813295430401,
	0.708731940200401,
	0.707648917255684,
	0.70656422914471,
	0.705477878419852,
	0.704389867637401,
	0.703300199357549,
	0.702208876144392,
	0.701115900565919,
	0.700021275194006,
	0.698925002604414,
	0.697827085376777,
	0.696727526094601,
	0.695626327345255,
	0.694523491719966,
	0.693419021813812,
	0.692312920225718,
	0.691205189558448,
	0.6900958324186,
	0.688984851416597,
	0.687872249166686,
	0.686758028286926,
	0.685642191399188,
	0.684524741129142,
	0.683405680106259,
	0.682285010963796,
	0.681162736338795,
	0.680038858872079,
	0.678913381208238,
	0.677786305995631,
	0.676657635886375,
	0.675527373536339,
	0.674395521605139,
	0.673262082756133,
	0.672127059656412,
	0.670990454976794,
	0.669852271391821,
	0.668712511579748,
	0.66757117822254,
	0.666428274005865,
	0.665283801619087,
	0.66413776375526,
	0.662990163111121,
	0.661841002387087,
	0.660690284287242,
	0.659538011519339,
	0.658384186794785,
	0.657228812828643,
	0.656071892339618,
	0.654913428050056,
	0.653753422685936,
	0.652591878976862,
	0.65142879965606,
	0.650264187460366,
	0.649098045130226,
	0.647930375409685,
	0.646761181046384,
	0.645590464791549,
	0.644418229399988,
	0.643244477630086,
	0.642069212243793,
	0.640892436006621,
	0.63971415168764,
	0.638534362059467,
	0.637353069898259,
	0.636170277983712,
	0.63498598909905,
	0.633800206031017,
	0.632612931569878,
	0.631424168509402,
	0.630233919646864,
	0.629042187783036,
	0.627848975722177,
	0.626654286272029,
	0.625458122243814,
	0.624260486452221,
	0.623061381715401,
	0.621860810854965,
	0.620658776695972,
	0.619455282066924,
	0.61825032979976,
	0.61704392272985,
	0.615836063695985,
	0.614626755540375,
	0.613416001108638,
	0.612203803249798,
	0.610990164816272,
	0.609775088663869,
	0.608558577651779,
	0.607340634642573,
	0.606121262502186,
	0.60490046409992,
	0.60367824230843,
	0.602454600003724,
	0.601229540065149,
	0.600003065375389,
	0.598775178820459,
	0.597545883289693,
	0.596315181675744,
	0.59508307687457,
	0.593849571785434,
	0.592614669310891,
	0.591378372356788,
	0.590140683832249,
	0.588901606649676,
	0.587661143724737,
	0.58641929797636,
	0.585176072326731,
	0.583931469701276,
	0.582685493028669,
	0.58143814524081,
	0.580189429272832,
	0.578939348063082,
	0.577687904553123,
	0.576435101687722,
	0.575180942414845,
	0.573925429685651,
	0.572668566454481,
	0.571410355678857,
	0.57015080031947,
	0.568889903340176,
	0.567627667707986,
	0.566364096393064,
	0.565099192368714,
	0.563832958611378,
	0.562565398100626,
	0.561296513819152,
	0.56002630875276,
	0.558754785890368,
	0.557481948223992,
	0.55620779874874,
	0.55493234046281,
	0.553655576367479,
	0.552377509467096,
	0.551098142769076,
	0.549817479283891,
	0.548535522025067,
	0.547252274009174,
	0.545967738255818,
	0.544681917787634,
	0.543394815630285,
	0.542106434812444,
	0.540816778365796,
	0.539525849325029,
	0.538233650727822,
	0.536940185614843,
	0.535645457029741,
	0.534349468019137,
	0.53305222163262,
	0.531753720922733,
	0.530453968944976,
	0.529152968757791,
	0.527850723422555,
	0.526547236003579,
	0.525242509568095,
	0.523936547186248,
	0.522629351931097,
	0.521320926878596,
	0.520011275107596,
	0.518700399699835,
	0.517388303739929,
	0.516074990315367,
	0.514760462516501,
	0.513444723436543,
	0.512127776171555,
	0.510809623820439,
	0.509490269484936,
	0.508169716269615,
	0.506847967281863,
	0.505525025631885,
	0.504200894432691,
	0.502875576800087,
	0.501549075852675,
	0.500221394711841,
	0.498892536501745,
	0.497562504349319,
	0.496231301384258,
	0.494898930739011,
	0.493565395548775,
	0.492230698951486,
	0.490894844087815,
	0.489557834101158,
	0.488219672137627,
	0.486880361346047,
	0.485539904877947,
	0.484198305887549,
	0.482855567531766,
	0.48151169297019,
	0.480166685365088,
	0.478820547881394,
	0.477473283686698,
	0.476124895951244,
	0.474775387847917,
	0.473424762552242,
	0.472073023242369,
	0.470720173099072,
	0.469366215305738,
	0.46801115304836,
	0.466654989515531,
	0.465297727898435,
	0.463939371390839,
	0.462579923189087,
	0.461219386492092,
	0.45985776450133,
	0.458495060420826,
	0.457131277457157,
	0.455766418819435,
	0.454400487719304,
	0.453033487370931,
	0.451665420991003,
	0.450296291798709,
	0.448926103015743,
	0.447554857866293,
	0.44618255957703,
	0.444809211377105,
	0.443434816498138,
	0.442059378174215,
	0.440682899641873,
	0.4393053841401,
	0.437926834910323,
	0.436547255196401,
	0.435166648244619,
	0.433785017303679,
	0.43240236562469,
	0.431018696461167,
	0.429634013069017,
	0.428248318706532,
	0.426861616634386,
	0.425473910115624,
	0.424085202415652,
	0.422695496802233,
	0.42130479654548,
	0.419913104917844,
	0.41852042519411,
	0.417126760651388,
	0.415732114569105,
	0.414336490228999,
	0.412939890915108,
	0.411542319913765,
	0.41014378051359,
	0.408744276005481,
	0.407343809682608,
	0.405942384840403,
	0.404540004776553,
	0.403136672790995,
	0.401732392185905,
	0.40032716626569,
	0.398920998336983,
	0.397513891708632,
	0.396105849691696,
	0.394696875599434,
	0.393286972747296,
	0.391876144452922,
	0.390464394036127,
	0.389051724818894,
	0.387638140125373,
	0.386223643281863,
	0.384808237616813,
	0.383391926460809,
	0.381974713146567,
	0.380556601008928,
	0.379137593384847,
	0.377717693613386,
	0.376296905035705,
	0.374875230995058,
	0.37345267483678,
	0.372029239908285,
	0.370604929559052,
	0.36917974714062,
	0.367753696006582,
	0.366326779512574,
	0.364899001016267,
	0.363470363877364,
	0.362040871457584,
	0.360610527120662,
	0.359179334232337,
	0.357747296160342,
	0.356314416274403,
	0.354880697946223,
	0.353446144549481,
	0.352010759459819,
	0.350574546054838,
	0.349137507714085,
	0.347699647819052,
	0.34626096975316,
	0.344821476901759,
	0.343381172652115,
	0.341940060393402,
	0.340498143516697,
	0.33905542541497,
	0.337611909483075,
	0.336167599117745,
	0.334722497717581,
	0.333276608683048,
	0.331829935416461,
	0.330382481321983,
	0.328934249805612,
	0.327485244275178,
	0.32603546814033,
	0.324584924812532,
	0.323133617705052,
	0.321681550232956,
	0.3202287258131,
	0.318775147864119,
	0.317320819806422,
	0.315865745062184,
	0.314409927055337,
	0.31295336921156,
	0.311496074958276,
	0.310038047724638,
	0.308579290941525,
	0.307119808041533,
	0.305659602458966,
	0.304198677629829,
	0.302737036991819,
	0.301274683984318,
	0.299811622048384,
	0.298347854626741,
	0.296883385163778,
	0.295418217105532,
	0.293952353899685,
	0.292485798995554,
	0.291018555844085,
	0.289550627897843,
	0.288082018611004,
	0.286612731439348,
	0.285142769840249,
	0.283672137272669,
	0.282200837197148,
	0.280728873075797,
	0.279256248372291,
	0.277782966551858,
	0.276309031081271,
	0.274834445428844,
	0.273359213064419,
	0.27188333745936,
	0.270406822086545,
	0.268929670420357,
	0.267451885936678,
	0.265973472112876,
	0.264494432427801,
	0.263014770361779,
	0.261534489396595,
	0.260053593015495,
	0.25857208470317,
	0.257089967945753,
	0.255607246230808,
	0.254123923047321,
	0.252640001885695,
	0.251155486237742,
	0.249670379596669,
	0.248184685457075,
	0.246698407314943,
	0.245211548667628,
	0.243724113013852,
	0.242236103853696,
	0.240747524688588,
	0.2392583790213,
	0.237768670355934,
	0.236278402197919,
	0.234787578054001,
	0.233296201432232,
	0.231804275841965,
	0.230311804793846,
	0.228818791799802,
	0.227325240373039,
	0.225831154028026,
	0.224336536280494,
	0.222841390647421,
	0.221345720647031,
	0.219849529798779,
	0.218352821623346,
	0.216855599642633,
	0.215357867379745,
	0.213859628358994,
	0.212360886105878,
	0.210861644147085,
	0.209361906010474,
	0.207861675225075,
	0.206360955321076,
	0.204859749829814,
	0.203358062283773,
	0.201855896216568,
	0.20035325516294,
	0.19885014265875,
	0.197346562240966,
	0.195842517447658,
	0.194338011817989,
	0.192833048892205,
	0.191327632211631,
	0.189821765318657,
	0.188315451756732,
	0.186808695070359,
	0.185301498805082,
	0.183793866507478,
	0.182285801725153,
	0.180777308006729,
	0.179268388901836,
	0.177759047961107,
	0.176249288736168,
	0.174739114779627,
	0.173228529645071,
	0.17171753688705,
	0.170206140061078,
	0.168694342723617,
	0.167182148432073,
	0.165669560744784,
	0.164156583221016,
	0.16264321942095,
	0.161129472905679,
	0.159615347237193,
	0.158100845978377,
	0.156585972692999,
	0.155070730945701,
	0.153555124301993,
	0.152039156328246,
	0.150522830591677,
	0.149006150660348,
	0.147489120103154,
	0.145971742489812,
	0.14445402139086,
	0.142935960377643,
	0.141417563022303,
	0.139898832897777,
	0.138379773577784,
	0.136860388636816,
	0.135340681650134,
	0.133820656193755,
	0.132300315844445,
	0.130779664179712,
	0.129258704777796,
	0.127737441217662,
	0.12621587707899,
	0.124694015942168,
	0.123171861388281,
	0.121649416999106,
	0.120126686357101,
	0.118603673045401,
	0.117080380647801,
	0.115556812748755,
	0.114032972933367,
	0.112508864787379,
	0.110984491897163,
	0.109459857849718,
	0.107934966232654,
	0.106409820634188,
	0.104884424643135,
	0.1033587818489,
	0.101832895841467,
	0.100306770211393,
	0.0987804085497995,
	0.0972538144483634,
	0.0957269914993072,
	0.094199943295393,
	0.0926726734299134,
	0.091145185496681,
	0.0896174830900232,
	0.0880895698047706,
	0.0865614492362511,
	0.0850331249802805,
	0.0835046006331525,
	0.0819758797916329,
	0.0804469660529502,
	0.0789178630147849,
	0.0773885742752649,
	0.0758591034329546,
	0.0743294540868457,
	0.0727996298363519,
	0.0712696342812965,
	0.0697394710219072,
	0.0682091436588065,
	0.0666786557930016,
	0.0651480110258787,
	0.0636172129591932,
	0.0620862651950601,
	0.0605551713359476,
	0.059023934984668,
	0.0574925597443675,
	0.0559610492185208,
	0.0544294070109192,
	0.0528976367256652,
	0.0513657419671628,
	0.0498337263401073,
	0.04830159344948,
	0.046769346900538,
	0.0452369902988046,
	0.0437045272500633,
	0.0421719613603481,
	0.0406392962359337,
	0.0391065354833301,
	0.0375736827092706,
	0.0360407415207061,
	0.034507715524796,
	0.0329746083288974,
	0.0314414235405602,
	0.0299081647675167,
	0.0283748356176721,
	0.0268414396990984,
	0.0253079806200247,
	0.0237744619888275,
	0.0222408874140252,
	0.020707260504266,
	0.0191735848683225,
	0.0176398641150823,
	0.0161061018535373,
	0.0145723016927789,
	0.0130384672419875,
	0.0115046021104227,
	0.00997070990741787,
	0.00843679424236992,
	0.00690285872472972,
	0.00536890696399659,
	0.00383494256970631,
	0.00230096915142573,
	0.000766990318742908,
	-0.000766990318742663,
	-0.00230096915142548,
	-0.00383494256970606,
	-0.00536890696399634,
	-0.00690285872472947,
	-0.00843679424236968,
	-0.00997070990741762,
	-0.0115046021104225,
	-0.0130384672419872,
	-0.0145723016927787,
	-0.0161061018535371,
	-0.017639864115082,
	-0.0191735848683223,
	-0.0207072605042657,
	-0.022240887414025,
	-0.0237744619888273,
	-0.0253079806200244,
	-0.0268414396990981,
	-0.0283748356176719,
	-0.0299081647675165,
	-0.0314414235405599,
	-0.0329746083288971,
	-0.0345077155247957,
	-0.0360407415207059,
	-0.0375736827092703,
	-0.0391065354833299,
	-0.0406392962359335,
	-0.0421719613603478,
	-0.043704527250063,
	-0.0452369902988043,
	-0.0467693469005378,
	-0.0483015934494798,
	-0.0498337263401071,
	-0.0513657419671625,
	-0.052897636725665,
	-0.054429407010919,
	-0.0559610492185206,
	-0.0574925597443673,
	-0.0590239349846678,
	-0.0605551713359474,
	-0.0620862651950598,
	-0.063617212959193,
	-0.0651480110258785,
	-0.0666786557930014,
	-0.0682091436588063,
	-0.069739471021907,
	-0.0712696342812962,
	-0.0727996298363517,
	-0.0743294540868455,
	-0.0758591034329543,
	-0.0773885742752646,
	-0.0789178630147847,
	-0.0804469660529499,
	-0.0819758797916327,
	-0.0835046006331522,
	-0.0850331249802802,
	-0.0865614492362508,
	-0.0880895698047703,
	-0.089617483090023,
	-0.0911451854966807,
	-0.0926726734299132,
	-0.0941999432953928,
	-0.0957269914993069,
	-0.0972538144483632,
	-0.0987804085497993,
	-0.100306770211393,
	-0.101832895841466,
	-0.103358781848899,
	-0.104884424643135,
	-0.106409820634188,
	-0.107934966232653,
	-0.109459857849718,
	-0.110984491897163,
	-0.112508864787378,
	-0.114032972933367,
	-0.115556812748755,
	-0.1170803806478,
	-0.118603673045401,
	-0.120126686357101,
	-0.121649416999105,
	-0.12317186138828,
	-0.124694015942167,
	-0.12621587707899,
	-0.127737441217662,
	-0.129258704777796,
	-0.130779664179712,
	-0.132300315844444,
	-0.133820656193755,
	-0.135340681650134,
	-0.136860388636816,
	-0.138379773577784,
	-0.139898832897777,
	-0.141417563022303,
	-0.142935960377643,
	-0.14445402139086,
	-0.145971742489812,
	-0.147489120103153,
	-0.149006150660348,
	-0.150522830591677,
	-0.152039156328246,
	-0.153555124301993,
	-0.1550707309457,
	-0.156585972692998,
	-0.158100845978377,
	-0.159615347237193,
	-0.161129472905678,
	-0.16264321942095,
	-0.164156583221016,
	-0.165669560744784,
	-0.167182148432073,
	-0.168694342723617,
	-0.170206140061078,
	-0.17171753688705,
	-0.17322852964507,
	-0.174739114779627,
	-0.176249288736168,
	-0.177759047961107,
	-0.179268388901835,
	-0.180777308006728,
	-0.182285801725153,
	-0.183793866507478,
	-0.185301498805082,
	-0.186808695070359,
	-0.188315451756732,
	-0.189821765318656,
	-0.191327632211631,
	-0.192833048892205,
	-0.194338011817989,
	-0.195842517447658,
	-0.197346562240966,
	-0.19885014265875,
	-0.20035325516294,
	-0.201855896216568,
	-0.203358062283773,
	-0.204859749829814,
	-0.206360955321075,
	-0.207861675225075,
	-0.209361906010474,
	-0.210861644147085,
	-0.212360886105878,
	-0.213859628358994,
	-0.215357867379745,
	-0.216855599642632,
	-0.218352821623346,
	-0.219849529798778,
	-0.221345720647031,
	-0.222841390647421,
	-0.224336536280493,
	-0.225831154028026,
	-0.227325240373039,
	-0.228818791799802,
	-0.230311804793845,
	-0.231804275841964,
	-0.233296201432231,
	-0.234787578054001,
	-0.236278402197919,
	-0.237768670355934,
	-0.2392583790213,
	-0.240747524688588,
	-0.242236103853696,
	-0.243724113013852,
	-0.245211548667627,
	-0.246698407314942,
	-0.248184685457074,
	-0.249670379596668,
	-0.251155486237742,
	-0.252640001885695,
	-0.25412392304732,
	-0.255607246230807,
	-0.257089967945753,
	-0.25857208470317,
	-0.260053593015495,
	-0.261534489396595,
	-0.263014770361779,
	-0.264494432427801,
	-0.265973472112875,
	-0.267451885936678,
	-0.268929670420357,
	-0.270406822086545,
	-0.27188333745936,
	-0.273359213064418,
	-0.274834445428844,
	-0.276309031081271,
	-0.277782966551857,
	-0.279256248372291,
	-0.280728873075797,
	-0.282200837197147,
	-0.283672137272668,
	-0.285142769840248,
	-0.286612731439348,
	-0.288082018611004,
	-0.289550627897843,
	-0.291018555844085,
	-0.292485798995554,
	-0.293952353899684,
	-0.295418217105532,
	-0.296883385163778,
	-0.298347854626741,
	-0.299811622048383,
	-0.301274683984318,
	-0.302737036991819,
	-0.304198677629829,
	-0.305659602458966,
	-0.307119808041533,
	-0.308579290941525,
	-0.310038047724638,
	-0.311496074958276,
	-0.31295336921156,
	-0.314409927055336,
	-0.315865745062184,
	-0.317320819806421,
	-0.318775147864118,
	-0.3202287258131,
	-0.321681550232956,
	-0.323133617705052,
	-0.324584924812532,
	-0.32603546814033,
	-0.327485244275178,
	-0.328934249805612,
	-0.330382481321983,
	-0.331829935416461,
	-0.333276608683048,
	-0.334722497717581,
	-0.336167599117744,
	-0.337611909483074,
	-0.339055425414969,
	-0.340498143516697,
	-0.341940060393402,
	-0.343381172652115,
	-0.344821476901759,
	-0.34626096975316,
	-0.347699647819051,
	-0.349137507714085,
	-0.350574546054837,
	-0.352010759459819,
	-0.35344614454948,
	-0.354880697946223,
	-0.356314416274402,
	-0.357747296160342,
	-0.359179334232336,
	-0.360610527120662,
	-0.362040871457584,
	-0.363470363877364,
	-0.364899001016267,
	-0.366326779512573,
	-0.367753696006582,
	-0.36917974714062,
	-0.370604929559051,
	-0.372029239908285,
	-0.37345267483678,
	-0.374875230995057,
	-0.376296905035704,
	-0.377717693613385,
	-0.379137593384847,
	-0.380556601008928,
	-0.381974713146567,
	-0.383391926460809,
	-0.384808237616813,
	-0.386223643281863,
	-0.387638140125373,
	-0.389051724818894,
	-0.390464394036126,
	-0.391876144452922,
	-0.393286972747296,
	-0.394696875599434,
	-0.396105849691696,
	-0.397513891708632,
	-0.398920998336983,
	-0.40032716626569,
	-0.401732392185905,
	-0.403136672790995,
	-0.404540004776553,
	-0.405942384840402,
	-0.407343809682608,
	-0.408744276005481,
	-0.41014378051359,
	-0.411542319913765,
	-0.412939890915108,
	-0.414336490228999,
	-0.415732114569105,
	-0.417126760651388,
	-0.41852042519411,
	-0.419913104917843,
	-0.42130479654548,
	-0.422695496802233,
	-0.424085202415651,
	-0.425473910115624,
	-0.426861616634386,
	-0.428248318706532,
	-0.429634013069016,
	-0.431018696461167,
	-0.43240236562469,
	-0.433785017303679,
	-0.435166648244619,
	-0.436547255196401,
	-0.437926834910323,
	-0.4393053841401,
	-0.440682899641873,
	-0.442059378174214,
	-0.443434816498138,
	-0.444809211377105,
	-0.44618255957703,
	-0.447554857866293,
	-0.448926103015743,
	-0.450296291798708,
	-0.451665420991002,
	-0.453033487370931,
	-0.454400487719303,
	-0.455766418819435,
	-0.457131277457157,
	-0.458495060420826,
	-0.459857764501329,
	-0.461219386492092,
	-0.462579923189087,
	-0.463939371390839,
	-0.465297727898434,
	-0.466654989515531,
	-0.468011153048359,
	-0.469366215305737,
	-0.470720173099072,
	-0.472073023242368,
	-0.473424762552241,
	-0.474775387847917,
	-0.476124895951243,
	-0.477473283686698,
	-0.478820547881394,
	-0.480166685365088,
	-0.48151169297019,
	-0.482855567531765,
	-0.484198305887549,
	-0.485539904877947,
	-0.486880361346047,
	-0.488219672137627,
	-0.489557834101157,
	-0.490894844087815,
	-0.492230698951486,
	-0.493565395548775,
	-0.494898930739011,
	-0.496231301384258,
	-0.497562504349319,
	-0.498892536501744,
	-0.500221394711841,
	-0.501549075852675,
	-0.502875576800087,
	-0.50420089443269,
	-0.505525025631885,
	-0.506847967281863,
	-0.508169716269615,
	-0.509490269484936,
	-0.510809623820439,
	-0.512127776171554,
	-0.513444723436543,
	-0.514760462516501,
	-0.516074990315366,
	-0.517388303739929,
	-0.518700399699835,
	-0.520011275107596,
	-0.521320926878595,
	-0.522629351931097,
	-0.523936547186248,
	-0.525242509568095,
	-0.526547236003579,
	-0.527850723422555,
	-0.529152968757791,
	-0.530453968944976,
	-0.531753720922733,
	-0.533052221632619,
	-0.534349468019137,
	-0.535645457029741,
	-0.536940185614843,
	-0.538233650727821,
	-0.539525849325029,
	-0.540816778365796,
	-0.542106434812444,
	-0.543394815630285,
	-0.544681917787634,
	-0.545967738255817,
	-0.547252274009174,
	-0.548535522025067,
	-0.549817479283891,
	-0.551098142769075,
	-0.552377509467096,
	-0.553655576367479,
	-0.55493234046281,
	-0.55620779874874,
	-0.557481948223991,
	-0.558754785890368,
	-0.56002630875276,
	-0.561296513819151,
	-0.562565398100626,
	-0.563832958611378,
	-0.565099192368714,
	-0.566364096393064,
	-0.567627667707986,
	-0.568889903340176,
	-0.57015080031947,
	-0.571410355678857,
	-0.572668566454481,
	-0.573925429685651,
	-0.575180942414845,
	-0.576435101687721,
	-0.577687904553123,
	-0.578939348063082,
	-0.580189429272831,
	-0.58143814524081,
	-0.582685493028668,
	-0.583931469701276,
	-0.58517607232673,
	-0.58641929797636,
	-0.587661143724736,
	-0.588901606649676,
	-0.590140683832249,
	-0.591378372356787,
	-0.592614669310891,
	-0.593849571785433,
	-0.59508307687457,
	-0.596315181675744,
	-0.597545883289693,
	-0.598775178820459,
	-0.600003065375389,
	-0.601229540065148,
	-0.602454600003724,
	-0.60367824230843,
	-0.60490046409992,
	-0.606121262502186,
	-0.607340634642573,
	-0.608558577651779,
	-0.609775088663868,
	-0.610990164816272,
	-0.612203803249798,
	-0.613416001108638,
	-0.614626755540375,
	-0.615836063695985,
	-0.617043922729849,
	-0.61825032979976,
	-0.619455282066924,
	-0.620658776695972,
	-0.621860810854965,
	-0.623061381715401,
	-0.62426048645222,
	-0.625458122243814,
	-0.626654286272029,
	-0.627848975722176,
	-0.629042187783036,
	-0.630233919646864,
	-0.631424168509402,
	-0.632612931569877,
	-0.633800206031017,
	-0.634985989099049,
	-0.636170277983712,
	-0.637353069898259,
	-0.638534362059467,
	-0.63971415168764,
	-0.640892436006621,
	-0.642069212243792,
	-0.643244477630086,
	-0.644418229399988,
	-0.645590464791549,
	-0.646761181046384,
	-0.647930375409685,
	-0.649098045130226,
	-0.650264187460366,
	-0.65142879965606,
	-0.652591878976862,
	-0.653753422685936,
	-0.654913428050056,
	-0.656071892339617,
	-0.657228812828642,
	-0.658384186794785,
	-0.659538011519338,
	-0.660690284287242,
	-0.661841002387087,
	-0.662990163111121,
	-0.66413776375526,
	-0.665283801619087,
	-0.666428274005865,
	-0.66757117822254,
	-0.668712511579748,
	-0.669852271391821,
	-0.670990454976794,
	-0.672127059656412,
	-0.673262082756133,
	-0.674395521605139,
	-0.675527373536338,
	-0.676657635886375,
	-0.677786305995631,
	-0.678913381208238,
	-0.680038858872079,
	-0.681162736338795,
	-0.682285010963795,
	-0.683405680106259,
	-0.684524741129142,
	-0.685642191399187,
	-0.686758028286926,
	-0.687872249166685,
	-0.688984851416597,
	-0.6900958324186,
	-0.691205189558448,
	-0.692312920225718,
	-0.693419021813812,
	-0.694523491719965,
	-0.695626327345255,
	-0.696727526094601,
	-0.697827085376777,
	-0.698925002604414,
	-0.700021275194006,
	-0.701115900565919,
	-0.702208876144392,
	-0.703300199357549,
	-0.7043898676374,
	-0.705477878419852,
	-0.706564229144709,
	-0.707648917255684,
	-0.7087319402004,
	-0.709813295430401,
	-0.710892980401152,
	-0.71197099257205,
	-0.713047329406429,
	-0.714121988371564,
	-0.71519496693868,
	-0.716266262582953,
	-0.717335872783521,
	-0.71840379502349,
	-0.719470026789933,
	-0.720534565573905,
	-0.721597408870444,
	-0.722658554178576,
	-0.723717999001323,
	-0.724775740845711,
	-0.72583177722277,
	-0.726886105647545,
	-0.727938723639099,
	-0.728989628720519,
	-0.730038818418926,
	-0.731086290265474,
	-0.732132041795361,
	-0.733176070547833,
	-0.734218374066188,
	-0.735258949897787,
	-0.736297795594053,
	-0.737334908710483,
	-0.738370286806648,
	-0.739403927446206,
	-0.740435828196898,
	-0.741465986630563,
	-0.742494400323139,
	-0.743521066854669,
	-0.744545983809307,
	-0.745569148775325,
	-0.746590559345117,
	-0.747610213115205,
	-0.748628107686245,
	-0.749644240663033,
	-0.750658609654511,
	-0.751671212273768,
	-0.752682046138055,
	-0.753691108868781,
	-0.754698398091524,
	-0.755703911436036,
	-0.756707646536246,
	-0.757709601030268,
	-0.758709772560407,
	-0.759708158773163,
	-0.760704757319236,
	-0.761699565853535,
	-0.762692582035177,
	-0.763683803527501,
	-0.764673227998067,
	-0.765660853118662,
	-0.76664667656531,
	-0.767630696018273,
	-0.768612909162058,
	-0.769593313685423,
	-0.77057190728138,
	-0.771548687647206,
	-0.772523652484441,
	-0.773496799498899,
	-0.77446812640067,
	-0.77543763090413,
	-0.77640531072794,
	-0.777371163595056,
	-0.778335187232733,
	-0.77929737937253,
	-0.780257737750316,
	-0.781216260106276,
	-0.782172944184912,
	-0.783127787735057,
	-0.784080788509869,
	-0.785031944266848,
	-0.78598125276783,
	-0.786928711779001,
	-0.7878743190709,
	-0.78881807241842,
	-0.789759969600819,
	-0.790700008401721,
	-0.791638186609125,
	-0.792574502015407,
	-0.793508952417326,
	-0.79444153561603,
	-0.795372249417061,
	-0.796301091630359,
	-0.797228060070268,
	-0.798153152555543,
	-0.799076366909352,
	-0.799997700959281,
	-0.800917152537344,
	-0.801834719479981,
	-0.802750399628068,
	-0.803664190826924,
	-0.804576090926307,
	-0.805486097780429,
	-0.806394209247956,
	-0.807300423192014,
	-0.808204737480195,
	-0.809107149984558,
	-0.810007658581641,
	-0.810906261152459,
	-0.811802955582515,
	-0.812697739761799,
	-0.813590611584798,
	-0.814481568950498,
	-0.815370609762391,
	-0.816257731928477,
	-0.817142933361273,
	-0.818026211977813,
	-0.818907565699659,
	-0.819786992452899,
	-0.820664490168157,
	-0.821540056780597,
	-0.822413690229926,
	-0.8232853884604,
	-0.824155149420828,
	-0.82502297106458,
	-0.825888851349587,
	-0.826752788238348,
	-0.827614779697938,
	-0.828474823700007,
	-0.829332918220788,
	-0.830189061241102,
	-0.831043250746362,
	-0.831895484726577,
	-0.832745761176359,
	-0.833594078094925,
	-0.834440433486103,
	-0.835284825358337,
	-0.836127251724692,
	-0.836967710602856,
	-0.837806200015151,
	-0.838642717988527,
	-0.839477262554578,
	-0.84030983174954,
	-0.841140423614297,
	-0.841969036194388,
	-0.842795667540004,
	-0.843620315706004,
	-0.84444297875191,
	-0.845263654741918,
	-0.846082341744897,
	-0.846899037834397,
	-0.847713741088654,
	-0.848526449590592,
	-0.84933716142783,
	-0.850145874692685,
	-0.850952587482175,
	-0.851757297898029,
	-0.852560004046684,
	-0.853360704039295,
	-0.854159395991739,
	-0.854956078024614,
	-0.855750748263254,
	-0.85654340483772,
	-0.857334045882815,
	-0.858122669538086,
	-0.858909273947823,
	-0.859693857261073,
	-0.860476417631632,
	-0.861256953218062,
	-0.862035462183687,
	-0.8628119426966,
	-0.863586392929668,
	-0.864358811060533,
	-0.865129195271623,
	-0.865897543750148,
	-0.866663854688111,
	-0.867428126282307,
	-0.868190356734331,
	-0.868950544250582,
	-0.869708687042265,
	-0.870464783325397,
	-0.871218831320811,
	-0.871970829254157,
	-0.872720775355914,
	-0.873468667861385,
	-0.874214505010706,
	-0.874958285048851,
	-0.875700006225634,
	-0.876439666795714,
	-0.877177265018596,
	-0.877912799158642,
	-0.878646267485068,
	-0.879377668271953,
	-0.88010699979824,
	-0.880834260347741,
	-0.881559448209143,
	-0.882282561676008,
	-0.883003599046781,
	-0.883722558624789,
	-0.884439438718253,
	-0.885154237640285,
	-0.885866953708892,
	-0.886577585246987,
	-0.887286130582383,
	-0.887992588047805,
	-0.888696955980892,
	-0.889399232724195,
	-0.890099416625192,
	-0.890797506036281,
	-0.891493499314791,
	-0.892187394822982,
	-0.892879190928051,
	-0.893568886002136,
	-0.894256478422316,
	-0.89494196657062,
	-0.89562534883403,
	-0.896306623604479,
	-0.896985789278864,
	-0.897662844259041,
	-0.898337786951834,
	-0.899010615769039,
	-0.899681329127423,
	-0.900349925448735,
	-0.901016403159702,
	-0.901680760692038,
	-0.902342996482444,
	-0.903003108972617,
	-0.903661096609248,
	-0.904316957844028,
	-0.904970691133653,
	-0.905622294939825,
	-0.906271767729257,
	-0.906919107973678,
	-0.907564314149832,
	-0.908207384739488,
	-0.908848318229439,
	-0.909487113111505,
	-0.910123767882542,
	-0.910758281044437,
	-0.911390651104122,
	-0.912020876573568,
	-0.912648955969794,
	-0.913274887814868,
	-0.913898670635911,
	-0.914520302965104,
	-0.915139783339685,
	-0.915757110301957,
	-0.916372282399289,
	-0.916985298184123,
	-0.917596156213973,
	-0.918204855051431,
	-0.91881139326417,
	-0.919415769424947,
	-0.920017982111606,
	-0.920618029907084,
	-0.921215911399408,
	-0.921811625181708,
	-0.92240516985221,
	-0.922996544014246,
	-0.923585746276257,
	-0.924172775251791,
	-0.924757629559514,
	-0.925340307823206,
	-0.92592080867177,
	-0.92649913073923,
	-0.92707527266474,
	-0.927649233092581,
	-0.928221010672169,
	-0.928790604058057,
	-0.929358011909935,
	-0.929923232892639,
	-0.930486265676149,
	-0.931047108935595,
	-0.931605761351258,
	-0.932162221608574,
	-0.93271648839814,
	-0.933268560415712,
	-0.933818436362211,
	-0.934366114943726,
	-0.934911594871516,
	-0.935454874862015,
	-0.935995953636831,
	-0.936534829922755,
	-0.937071502451759,
	-0.937605969961,
	-0.938138231192824,
	-0.93866828489477,
	-0.939196129819569,
	-0.939721764725153,
	-0.940245188374651,
	-0.940766399536396,
	-0.941285396983929,
	-0.941802179495997,
	-0.942316745856563,
	-0.942829094854802,
	-0.943339225285107,
	-0.943847135947093,
	-0.944352825645594,
	-0.944856293190677,
	-0.945357537397632,
	-0.945856557086984,
	-0.94635335108449,
	-0.946847918221148,
	-0.947340257333192,
	-0.947830367262101,
	-0.948318246854599,
	-0.948803894962658,
	-0.949287310443502,
	-0.949768492159607,
	-0.950247438978705,
	-0.950724149773789,
	-0.951198623423113,
	-0.951670858810194,
	-0.952140854823816,
	-0.952608610358033,
	-0.953074124312172,
	-0.953537395590833,
	-0.953998423103894,
	-0.954457205766513,
	-0.95491374249913,
	-0.95536803222747,
	-0.955820073882545,
	-0.956269866400658,
	-0.956717408723403,
	-0.95716269979767,
	-0.957605738575646,
	-0.958046524014818,
	-0.958485055077976,
	-0.958921330733213,
	-0.959355349953931,
	-0.95978711171884,
	-0.960216615011963,
	-0.960643858822638,
	-0.961068842145519,
	-0.961491563980579,
	-0.961912023333112,
	-0.962330219213737,
	-0.962746150638399,
	-0.963159816628371,
	-0.963571216210257,
	-0.963980348415994,
	-0.964387212282854,
	-0.964791806853448,
	-0.965194131175725,
	-0.965594184302977,
	-0.96599196529384,
	-0.966387473212299,
	-0.966780707127683,
	-0.967171666114676,
	-0.967560349253314,
	-0.967946755628988,
	-0.968330884332445,
	-0.968712734459795,
	-0.969092305112506,
	-0.969469595397413,
	-0.969844604426715,
	-0.970217331317979,
	-0.970587775194144,
	-0.970955935183518,
	-0.971321810419786,
	-0.971685400042008,
	-0.972046703194623,
	-0.97240571902745,
	-0.972762446695688,
	-0.973116885359925,
	-0.973469034186131,
	-0.973818892345666,
	-0.97416645901528,
	-0.974511733377116,
	-0.974854714618708,
	-0.97519540193299,
	-0.975533794518291,
	-0.975869891578341,
	-0.97620369232227,
	-0.976535195964614,
	-0.976864401725312,
	-0.977191308829712,
	-0.977515916508569,
	-0.97783822399805,
	-0.978158230539735,
	-0.978475935380617,
	-0.978791337773105,
	-0.979104436975029,
	-0.979415232249635,
	-0.979723722865591,
	-0.98002990809699,
	-0.980333787223348,
	-0.980635359529608,
	-0.980934624306142,
	-0.98123158084875,
	-0.981526228458665,
	-0.981818566442552,
	-0.982108594112513,
	-0.982396310786085,
	-0.982681715786241,
	-0.982964808441396,
	-0.983245588085407,
	-0.983524054057571,
	-0.983800205702631,
	-0.984074042370776,
	-0.984345563417642,
	-0.984614768204312,
	-0.984881656097323,
	-0.985146226468662,
	-0.985408478695768,
	-0.985668412161537,
	-0.985926026254321,
	-0.986181320367928,
	-0.986434293901627,
	-0.986684946260147,
	-0.986933276853678,
	-0.987179285097874,
	-0.987422970413855,
	-0.987664332228206,
	-0.987903369972978,
	-0.988140083085692,
	-0.988374471009341,
	-0.988606533192386,
	-0.988836269088763,
	-0.989063678157881,
	-0.989288759864625,
	-0.989511513679355,
	-0.989731939077911,
	-0.989950035541609,
	-0.990165802557248,
	-0.990379239617108,
	-0.99059034621895,
	-0.99079912186602,
	-0.991005566067049,
	-0.991209678336254,
	-0.991411458193339,
	-0.991610905163495,
	-0.991808018777406,
	-0.992002798571245,
	-0.992195244086674,
	-0.992385354870852,
	-0.992573130476429,
	-0.992758570461551,
	-0.99294167438986,
	-0.993122441830496,
	-0.993300872358093,
	-0.993476965552789,
	-0.993650721000219,
	-0.99382213829152,
	-0.993991217023329,
	-0.99415795679779,
	-0.994322357222546,
	-0.994484417910747,
	-0.994644138481051,
	-0.994801518557617,
	-0.994956557770116,
	-0.995109255753726,
	-0.995259612149133,
	-0.995407626602535,
	-0.995553298765638,
	-0.995696628295663,
	-0.995837614855342,
	-0.995976258112918,
	-0.996112557742151,
	-0.996246513422315,
	-0.9963781248382,
	-0.996507391680111,
	-0.99663431364387,
	-0.996758890430818,
	-0.996881121747814,
	-0.997001007307235,
	-0.99711854682698,
	-0.997233740030466,
	-0.997346586646633,
	-0.997457086409942,
	-0.997565239060376,
	-0.997671044343441,
	-0.997774502010168,
	-0.99787561181711,
	-0.997974373526347,
	-0.998070786905482,
	-0.998164851727646,
	-0.998256567771495,
	-0.998345934821212,
	-0.998432952666508,
	-0.998517621102622,
	-0.99859993993032,
	-0.998679908955899,
	-0.998757527991183,
	-0.998832796853528,
	-0.998905715365818,
	-0.99897628335647,
	-0.999044500659429,
	-0.999110367114175,
	-0.999173882565716,
	-0.999235046864596,
	-0.999293859866888,
	-0.999350321434199,
	-0.999404431433671,
	-0.999456189737977,
	-0.999505596225325,
	-0.999552650779457,
	-0.999597353289648,
	-0.99963970365071,
	-0.999679701762988,
	-0.999717347532362,
	-0.999752640870249,
	-0.999785581693599,
	-0.9998161699249,
	-0.999844405492175,
	-0.999870288328983,
	-0.999893818374418,
	-0.999914995573113,
	-0.999933819875236,
	-0.99995029123649,
	-0.999964409618118,
	-0.999976174986898,
	-0.999985587315143,
	-0.999992646580707,
	-0.999997352766978,
	-0.999999705862882,
	-0.999999705862882,
	-0.999997352766978,
	-0.999992646580707,
	-0.999985587315143,
	-0.999976174986898,
	-0.999964409618118,
	-0.99995029123649,
	-0.999933819875236,
	-0.999914995573114,
	-0.999893818374418,
	-0.999870288328983,
	-0.999844405492175,
	-0.9998161699249,
	-0.999785581693599,
	-0.999752640870249,
	-0.999717347532362,
	-0.999679701762988,
	-0.99963970365071,
	-0.999597353289648,
	-0.999552650779457,
	-0.999505596225325,
	-0.999456189737977,
	-0.999404431433671,
	-0.999350321434199,
	-0.999293859866888,
	-0.999235046864596,
	-0.999173882565716,
	-0.999110367114175,
	-0.999044500659429,
	-0.99897628335647,
	-0.998905715365818,
	-0.998832796853528,
	-0.998757527991183,
	-0.998679908955899,
	-0.99859993993032,
	-0.998517621102622,
	-0.998432952666509,
	-0.998345934821212,
	-0.998256567771495,
	-0.998164851727646,
	-0.998070786905482,
	-0.997974373526347,
	-0.99787561181711,
	-0.997774502010168,
	-0.997671044343441,
	-0.997565239060376,
	-0.997457086409942,
	-0.997346586646633,
	-0.997233740030466,
	-0.99711854682698,
	-0.997001007307235,
	-0.996881121747814,
	-0.996758890430818,
	-0.99663431364387,
	-0.996507391680111,
	-0.9963781248382,
	-0.996246513422316,
	-0.996112557742151,
	-0.995976258112918,
	-0.995837614855342,
	-0.995696628295664,
	-0.995553298765639,
	-0.995407626602535,
	-0.995259612149133,
	-0.995109255753726,
	-0.994956557770116,
	-0.994801518557617,
	-0.994644138481051,
	-0.994484417910748,
	-0.994322357222546,
	-0.99415795679779,
	-0.993991217023329,
	-0.99382213829152,
	-0.993650721000219,
	-0.993476965552789,
	-0.993300872358093,
	-0.993122441830496,
	-0.992941674389861,
	-0.992758570461551,
	-0.992573130476429,
	-0.992385354870852,
	-0.992195244086674,
	-0.992002798571245,
	-0.991808018777407,
	-0.991610905163495,
	-0.991411458193339,
	-0.991209678336254,
	-0.991005566067049,
	-0.99079912186602,
	-0.99059034621895,
	-0.990379239617108,
	-0.990165802557249,
	-0.989950035541609,
	-0.989731939077911,
	-0.989511513679355,
	-0.989288759864625,
	-0.989063678157882,
	-0.988836269088764,
	-0.988606533192387,
	-0.988374471009341,
	-0.988140083085693,
	-0.987903369972978,
	-0.987664332228206,
	-0.987422970413856,
	-0.987179285097874,
	-0.986933276853678,
	-0.986684946260147,
	-0.986434293901627,
	-0.986181320367928,
	-0.985926026254321,
	-0.985668412161538,
	-0.985408478695769,
	-0.985146226468662,
	-0.984881656097324,
	-0.984614768204313,
	-0.984345563417642,
	-0.984074042370777,
	-0.983800205702632,
	-0.983524054057571,
	-0.983245588085407,
	-0.982964808441397,
	-0.982681715786241,
	-0.982396310786085,
	-0.982108594112514,
	-0.981818566442553,
	-0.981526228458665,
	-0.98123158084875,
	-0.980934624306142,
	-0.980635359529608,
	-0.980333787223348,
	-0.98002990809699,
	-0.979723722865591,
	-0.979415232249635,
	-0.979104436975029,
	-0.978791337773106,
	-0.978475935380617,
	-0.978158230539735,
	-0.977838223998051,
	-0.977515916508569,
	-0.977191308829712,
	-0.976864401725313,
	-0.976535195964615,
	-0.976203692322271,
	-0.975869891578341,
	-0.975533794518291,
	-0.975195401932991,
	-0.974854714618709,
	-0.974511733377116,
	-0.974166459015281,
	-0.973818892345666,
	-0.973469034186131,
	-0.973116885359925,
	-0.972762446695689,
	-0.97240571902745,
	-0.972046703194624,
	-0.971685400042009,
	-0.971321810419786,
	-0.970955935183518,
	-0.970587775194144,
	-0.970217331317979,
	-0.969844604426715,
	-0.969469595397413,
	-0.969092305112506,
	-0.968712734459795,
	-0.968330884332445,
	-0.967946755628988,
	-0.967560349253314,
	-0.967171666114677,
	-0.966780707127684,
	-0.966387473212299,
	-0.965991965293841,
	-0.965594184302977,
	-0.965194131175725,
	-0.964791806853448,
	-0.964387212282855,
	-0.963980348415994,
	-0.963571216210257,
	-0.963159816628371,
	-0.9627461506384,
	-0.962330219213738,
	-0.961912023333112,
	-0.961491563980579,
	-0.961068842145519,
	-0.960643858822639,
	-0.960216615011964,
	-0.95978711171884,
	-0.959355349953931,
	-0.958921330733213,
	-0.958485055077976,
	-0.958046524014819,
	-0.957605738575647,
	-0.95716269979767,
	-0.956717408723403,
	-0.956269866400658,
	-0.955820073882546,
	-0.95536803222747,
	-0.954913742499131,
	-0.954457205766514,
	-0.953998423103895,
	-0.953537395590833,
	-0.953074124312172,
	-0.952608610358034,
	-0.952140854823816,
	-0.951670858810194,
	-0.951198623423113,
	-0.95072414977379,
	-0.950247438978706,
	-0.949768492159607,
	-0.949287310443502,
	-0.948803894962659,
	-0.948318246854599,
	-0.947830367262101,
	-0.947340257333192,
	-0.946847918221148,
	-0.946353351084491,
	-0.945856557086984,
	-0.945357537397633,
	-0.944856293190677,
	-0.944352825645595,
	-0.943847135947093,
	-0.943339225285108,
	-0.942829094854803,
	-0.942316745856564,
	-0.941802179495998,
	-0.941285396983929,
	-0.940766399536396,
	-0.940245188374651,
	-0.939721764725153,
	-0.93919612981957,
	-0.93866828489477,
	-0.938138231192825,
	-0.937605969961,
	-0.937071502451759,
	-0.936534829922756,
	-0.935995953636832,
	-0.935454874862015,
	-0.934911594871516,
	-0.934366114943726,
	-0.933818436362211,
	-0.933268560415712,
	-0.932716488398141,
	-0.932162221608575,
	-0.931605761351258,
	-0.931047108935595,
	-0.93048626567615,
	-0.92992323289264,
	-0.929358011909936,
	-0.928790604058057,
	-0.92822101067217,
	-0.927649233092581,
	-0.927075272664741,
	-0.926499130739231,
	-0.92592080867177,
	-0.925340307823207,
	-0.924757629559514,
	-0.924172775251792,
	-0.923585746276257,
	-0.922996544014247,
	-0.92240516985221,
	-0.921811625181708,
	-0.921215911399409,
	-0.920618029907084,
	-0.920017982111607,
	-0.919415769424947,
	-0.91881139326417,
	-0.918204855051431,
	-0.917596156213973,
	-0.916985298184123,
	-0.916372282399289,
	-0.915757110301957,
	-0.915139783339685,
	-0.914520302965105,
	-0.913898670635912,
	-0.913274887814868,
	-0.912648955969794,
	-0.912020876573569,
	-0.911390651104123,
	-0.910758281044438,
	-0.910123767882542,
	-0.909487113111506,
	-0.908848318229439,
	-0.908207384739489,
	-0.907564314149833,
	-0.906919107973678,
	-0.906271767729258,
	-0.905622294939826,
	-0.904970691133653,
	-0.904316957844029,
	-0.903661096609248,
	-0.903003108972618,
	-0.902342996482445,
	-0.901680760692038,
	-0.901016403159703,
	-0.900349925448736,
	-0.899681329127424,
	-0.89901061576904,
	-0.898337786951835,
	-0.897662844259041,
	-0.896985789278864,
	-0.89630662360448,
	-0.895625348834031,
	-0.894941966570621,
	-0.894256478422316,
	-0.893568886002136,
	-0.892879190928052,
	-0.892187394822983,
	-0.891493499314792,
	-0.890797506036282,
	-0.890099416625193,
	-0.889399232724196,
	-0.888696955980892,
	-0.887992588047806,
	-0.887286130582384,
	-0.886577585246987,
	-0.885866953708893,
	-0.885154237640285,
	-0.884439438718254,
	-0.88372255862479,
	-0.883003599046781,
	-0.882282561676009,
	-0.881559448209144,
	-0.880834260347743,
	-0.880106999798241,
	-0.879377668271954,
	-0.878646267485068,
	-0.877912799158642,
	-0.877177265018597,
	-0.876439666795714,
	-0.875700006225635,
	-0.874958285048852,
	-0.874214505010707,
	-0.873468667861385,
	-0.872720775355914,
	-0.871970829254158,
	-0.871218831320811,
	-0.870464783325398,
	-0.869708687042266,
	-0.868950544250583,
	-0.868190356734332,
	-0.867428126282307,
	-0.866663854688111,
	-0.865897543750149,
	-0.865129195271624,
	-0.864358811060535,
	-0.863586392929669,
	-0.862811942696601,
	-0.862035462183688,
	-0.861256953218063,
	-0.860476417631633,
	-0.859693857261073,
	-0.858909273947824,
	-0.858122669538087,
	-0.857334045882816,
	-0.85654340483772,
	-0.855750748263254,
	-0.854956078024615,
	-0.854159395991739,
	-0.853360704039296,
	-0.852560004046684,
	-0.851757297898029,
	-0.850952587482176,
	-0.850145874692686,
	-0.849337161427831,
	-0.848526449590593,
	-0.847713741088655,
	-0.846899037834398,
	-0.846082341744897,
	-0.845263654741919,
	-0.844442978751911,
	-0.843620315706004,
	-0.842795667540005,
	-0.841969036194388,
	-0.841140423614299,
	-0.840309831749541,
	-0.839477262554579,
	-0.838642717988528,
	-0.837806200015151,
	-0.836967710602858,
	-0.836127251724693,
	-0.835284825358338,
	-0.834440433486103,
	-0.833594078094925,
	-0.83274576117636,
	-0.831895484726578,
	-0.831043250746363,
	-0.830189061241103,
	-0.829332918220788,
	-0.828474823700008,
	-0.827614779697939,
	-0.826752788238349,
	-0.825888851349587,
	-0.825022971064581,
	-0.824155149420829,
	-0.823285388460401,
	-0.822413690229927,
	-0.821540056780598,
	-0.820664490168158,
	-0.819786992452899,
	-0.818907565699659,
	-0.818026211977814,
	-0.817142933361274,
	-0.816257731928478,
	-0.815370609762392,
	-0.814481568950499,
	-0.813590611584799,
	-0.8126977397618,
	-0.811802955582516,
	-0.81090626115246,
	-0.810007658581641,
	-0.809107149984559,
	-0.808204737480195,
	-0.807300423192015,
	-0.806394209247957,
	-0.805486097780429,
	-0.804576090926307,
	-0.803664190826924,
	-0.80275039962807,
	-0.801834719479982,
	-0.800917152537345,
	-0.799997700959282,
	-0.799076366909353,
	-0.798153152555544,
	-0.797228060070269,
	-0.79630109163036,
	-0.795372249417062,
	-0.794441535616031,
	-0.793508952417327,
	-0.792574502015408,
	-0.791638186609126,
	-0.790700008401722,
	-0.789759969600819,
	-0.788818072418421,
	-0.787874319070901,
	-0.786928711779002,
	-0.785981252767831,
	-0.785031944266848,
	-0.78408078850987,
	-0.783127787735057,
	-0.782172944184914,
	-0.781216260106277,
	-0.780257737750317,
	-0.779297379372531,
	-0.778335187232733,
	-0.777371163595057,
	-0.776405310727941,
	-0.775437630904131,
	-0.774468126400671,
	-0.773496799498899,
	-0.772523652484442,
	-0.771548687647207,
	-0.770571907281381,
	-0.769593313685423,
	-0.768612909162059,
	-0.767630696018274,
	-0.766646676565311,
	-0.765660853118663,
	-0.764673227998068,
	-0.763683803527502,
	-0.762692582035178,
	-0.761699565853535,
	-0.760704757319238,
	-0.759708158773164,
	-0.758709772560408,
	-0.757709601030268,
	-0.756707646536246,
	-0.755703911436037,
	-0.754698398091525,
	-0.753691108868782,
	-0.752682046138056,
	-0.751671212273769,
	-0.750658609654511,
	-0.749644240663034,
	-0.748628107686246,
	-0.747610213115206,
	-0.746590559345118,
	-0.745569148775326,
	-0.744545983809308,
	-0.74352106685467,
	-0.74249440032314,
	-0.741465986630564,
	-0.740435828196898,
	-0.739403927446206,
	-0.738370286806649,
	-0.737334908710483,
	-0.736297795594054,
	-0.735258949897787,
	-0.734218374066189,
	-0.733176070547834,
	-0.732132041795362,
	-0.731086290265475,
	-0.730038818418927,
	-0.72898962872052,
	-0.727938723639099,
	-0.726886105647546,
	-0.725831777222771,
	-0.724775740845712,
	-0.723717999001324,
	-0.722658554178576,
	-0.721597408870444,
	-0.720534565573906,
	-0.719470026789934,
	-0.71840379502349,
	-0.717335872783522,
	-0.716266262582953,
	-0.715194966938681,
	-0.714121988371565,
	-0.71304732940643,
	-0.71197099257205,
	-0.710892980401152,
	-0.709813295430402,
	-0.708731940200401,
	-0.707648917255685,
	-0.70656422914471,
	-0.705477878419852,
	-0.704389867637401,
	-0.703300199357549,
	-0.702208876144392,
	-0.701115900565919,
	-0.700021275194007,
	-0.698925002604415,
	-0.697827085376778,
	-0.696727526094602,
	-0.695626327345255,
	-0.694523491719966,
	-0.693419021813812,
	-0.692312920225718,
	-0.691205189558449,
	-0.690095832418601,
	-0.688984851416597,
	-0.687872249166686,
	-0.686758028286926,
	-0.685642191399188,
	-0.684524741129143,
	-0.683405680106259,
	-0.682285010963796,
	-0.681162736338796,
	-0.68003885887208,
	-0.678913381208239,
	-0.677786305995632,
	-0.676657635886375,
	-0.675527373536339,
	-0.67439552160514,
	-0.673262082756134,
	-0.672127059656412,
	-0.670990454976795,
	-0.669852271391821,
	-0.668712511579748,
	-0.667571178222541,
	-0.666428274005866,
	-0.665283801619088,
	-0.66413776375526,
	-0.662990163111122,
	-0.661841002387087,
	-0.660690284287243,
	-0.659538011519339,
	-0.658384186794786,
	-0.657228812828643,
	-0.656071892339618,
	-0.654913428050057,
	-0.653753422685937,
	-0.652591878976863,
	-0.65142879965606,
	-0.650264187460366,
	-0.649098045130227,
	-0.647930375409686,
	-0.646761181046385,
	-0.645590464791549,
	-0.644418229399989,
	-0.643244477630086,
	-0.642069212243793,
	-0.640892436006622,
	-0.639714151687641,
	-0.638534362059467,
	-0.63735306989826,
	-0.636170277983712,
	-0.63498598909905,
	-0.633800206031018,
	-0.632612931569878,
	-0.631424168509402,
	-0.630233919646865,
	-0.629042187783037,
	-0.627848975722177,
	-0.62665428627203,
	-0.625458122243815,
	-0.624260486452221,
	-0.623061381715402,
	-0.621860810854966,
	-0.620658776695973,
	-0.619455282066925,
	-0.618250329799761,
	-0.61704392272985,
	-0.615836063695985,
	-0.614626755540376,
	-0.613416001108639,
	-0.612203803249799,
	-0.610990164816272,
	-0.609775088663869,
	-0.60855857765178,
	-0.607340634642574,
	-0.606121262502187,
	-0.60490046409992,
	-0.603678242308431,
	-0.602454600003725,
	-0.601229540065149,
	-0.60000306537539,
	-0.598775178820459,
	-0.597545883289694,
	-0.596315181675745,
	-0.595083076874571,
	-0.593849571785434,
	-0.592614669310892,
	-0.591378372356788,
	-0.590140683832249,
	-0.588901606649676,
	-0.587661143724738,
	-0.586419297976361,
	-0.585176072326731,
	-0.583931469701277,
	-0.582685493028669,
	-0.581438145240811,
	-0.580189429272832,
	-0.578939348063082,
	-0.577687904553123,
	-0.576435101687722,
	-0.575180942414846,
	-0.573925429685652,
	-0.572668566454482,
	-0.571410355678858,
	-0.570150800319471,
	-0.568889903340176,
	-0.567627667707987,
	-0.566364096393065,
	-0.565099192368715,
	-0.563832958611379,
	-0.562565398100627,
	-0.561296513819152,
	-0.560026308752761,
	-0.558754785890369,
	-0.557481948223992,
	-0.55620779874874,
	-0.554932340462811,
	-0.55365557636748,
	-0.552377509467097,
	-0.551098142769076,
	-0.549817479283891,
	-0.548535522025068,
	-0.547252274009175,
	-0.545967738255818,
	-0.544681917787635,
	-0.543394815630285,
	-0.542106434812444,
	-0.540816778365797,
	-0.53952584932503,
	-0.538233650727822,
	-0.536940185614844,
	-0.535645457029742,
	-0.534349468019138,
	-0.53305222163262,
	-0.531753720922734,
	-0.530453968944977,
	-0.529152968757791,
	-0.527850723422556,
	-0.52654723600358,
	-0.525242509568096,
	-0.523936547186249,
	-0.522629351931097,
	-0.521320926878596,
	-0.520011275107596,
	-0.518700399699836,
	-0.51738830373993,
	-0.516074990315367,
	-0.514760462516502,
	-0.513444723436544,
	-0.512127776171555,
	-0.51080962382044,
	-0.509490269484937,
	-0.508169716269615,
	-0.506847967281864,
	-0.505525025631886,
	-0.504200894432691,
	-0.502875576800088,
	-0.501549075852676,
	-0.500221394711841,
	-0.498892536501745,
	-0.497562504349319,
	-0.496231301384259,
	-0.494898930739012,
	-0.493565395548775,
	-0.492230698951487,
	-0.490894844087816,
	-0.489557834101158,
	-0.488219672137628,
	-0.486880361346048,
	-0.485539904877948,
	-0.48419830588755,
	-0.482855567531766,
	-0.481511692970191,
	-0.480166685365089,
	-0.478820547881395,
	-0.477473283686699,
	-0.476124895951244,
	-0.474775387847917,
	-0.473424762552242,
	-0.472073023242369,
	-0.470720173099072,
	-0.469366215305738,
	-0.46801115304836,
	-0.466654989515532,
	-0.465297727898435,
	-0.463939371390839,
	-0.462579923189087,
	-0.461219386492093,
	-0.459857764501331,
	-0.458495060420827,
	-0.457131277457158,
	-0.455766418819435,
	-0.454400487719304,
	-0.453033487370932,
	-0.451665420991003,
	-0.45029629179871,
	-0.448926103015744,
	-0.447554857866294,
	-0.44618255957703,
	-0.444809211377105,
	-0.443434816498139,
	-0.442059378174216,
	-0.440682899641874,
	-0.4393053841401,
	-0.437926834910323,
	-0.436547255196402,
	-0.43516664824462,
	-0.433785017303679,
	-0.432402365624691,
	-0.431018696461167,
	-0.429634013069017,
	-0.428248318706533,
	-0.426861616634387,
	-0.425473910115625,
	-0.424085202415652,
	-0.422695496802233,
	-0.421304796545481,
	-0.419913104917845,
	-0.41852042519411,
	-0.417126760651388,
	-0.415732114569106,
	-0.414336490228999,
	-0.412939890915109,
	-0.411542319913766,
	-0.410143780513591,
	-0.408744276005482,
	-0.407343809682608,
	-0.405942384840404,
	-0.404540004776554,
	-0.403136672790996,
	-0.401732392185906,
	-0.400327166265691,
	-0.398920998336984,
	-0.397513891708633,
	-0.396105849691697,
	-0.394696875599434,
	-0.393286972747297,
	-0.391876144452923,
	-0.390464394036128,
	-0.389051724818895,
	-0.387638140125373,
	-0.386223643281864,
	-0.384808237616813,
	-0.383391926460809,
	-0.381974713146568,
	-0.380556601008929,
	-0.379137593384848,
	-0.377717693613386,
	-0.376296905035705,
	-0.374875230995059,
	-0.373452674836781,
	-0.372029239908286,
	-0.370604929559052,
	-0.36917974714062,
	-0.367753696006583,
	-0.366326779512575,
	-0.364899001016268,
	-0.363470363877364,
	-0.362040871457585,
	-0.360610527120663,
	-0.359179334232338,
	-0.357747296160343,
	-0.356314416274403,
	-0.354880697946223,
	-0.353446144549481,
	-0.352010759459819,
	-0.350574546054839,
	-0.349137507714086,
	-0.347699647819052,
	-0.346260969753161,
	-0.34482147690176,
	-0.343381172652116,
	-0.341940060393403,
	-0.340498143516698,
	-0.33905542541497,
	-0.337611909483075,
	-0.336167599117746,
	-0.334722497717582,
	-0.333276608683049,
	-0.331829935416462,
	-0.330382481321983,
	-0.328934249805613,
	-0.327485244275179,
	-0.326035468140331,
	-0.324584924812533,
	-0.323133617705053,
	-0.321681550232957,
	-0.3202287258131,
	-0.31877514786412,
	-0.317320819806423,
	-0.315865745062185,
	-0.314409927055337,
	-0.312953369211561,
	-0.311496074958277,
	-0.310038047724639,
	-0.308579290941526,
	-0.307119808041534,
	-0.305659602458967,
	-0.30419867762983,
	-0.30273703699182,
	-0.301274683984319,
	-0.299811622048384,
	-0.298347854626742,
	-0.296883385163779,
	-0.295418217105533,
	-0.293952353899686,
	-0.292485798995555,
	-0.291018555844086,
	-0.289550627897844,
	-0.288082018611004,
	-0.286612731439349,
	-0.28514276984025,
	-0.283672137272669,
	-0.282200837197148,
	-0.280728873075798,
	-0.279256248372292,
	-0.277782966551859,
	-0.276309031081272,
	-0.274834445428845,
	-0.273359213064419,
	-0.271883337459361,
	-0.270406822086546,
	-0.268929670420358,
	-0.267451885936678,
	-0.265973472112876,
	-0.264494432427802,
	-0.26301477036178,
	-0.261534489396596,
	-0.260053593015496,
	-0.258572084703171,
	-0.257089967945754,
	-0.255607246230808,
	-0.254123923047322,
	-0.252640001885696,
	-0.251155486237743,
	-0.249670379596669,
	-0.248184685457075,
	-0.246698407314944,
	-0.245211548667629,
	-0.243724113013853,
	-0.242236103853697,
	-0.240747524688589,
	-0.2392583790213,
	-0.237768670355935,
	-0.23627840219792,
	-0.234787578054002,
	-0.233296201432232,
	-0.231804275841965,
	-0.230311804793847,
	-0.228818791799803,
	-0.22732524037304,
	-0.225831154028027,
	-0.224336536280494,
	-0.222841390647421,
	-0.221345720647032,
	-0.21984952979878,
	-0.218352821623347,
	-0.216855599642633,
	-0.215357867379746,
	-0.213859628358995,
	-0.212360886105879,
	-0.210861644147086,
	-0.209361906010475,
	-0.207861675225076,
	-0.206360955321076,
	-0.204859749829815,
	-0.203358062283774,
	-0.201855896216569,
	-0.200353255162941,
	-0.198850142658751,
	-0.197346562240967,
	-0.195842517447659,
	-0.194338011817989,
	-0.192833048892206,
	-0.191327632211631,
	-0.189821765318657,
	-0.188315451756733,
	-0.18680869507036,
	-0.185301498805083,
	-0.183793866507479,
	-0.182285801725154,
	-0.18077730800673,
	-0.179268388901837,
	-0.177759047961108,
	-0.176249288736169,
	-0.174739114779628,
	-0.173228529645071,
	-0.171717536887051,
	-0.170206140061079,
	-0.168694342723618,
	-0.167182148432074,
	-0.165669560744785,
	-0.164156583221017,
	-0.162643219420951,
	-0.16112947290568,
	-0.159615347237194,
	-0.158100845978378,
	-0.156585972692999,
	-0.155070730945702,
	-0.153555124301994,
	-0.152039156328247,
	-0.150522830591678,
	-0.149006150660349,
	-0.147489120103155,
	-0.145971742489813,
	-0.144454021390861,
	-0.142935960377643,
	-0.141417563022304,
	-0.139898832897778,
	-0.138379773577785,
	-0.136860388636817,
	-0.135340681650135,
	-0.133820656193755,
	-0.132300315844445,
	-0.130779664179713,
	-0.129258704777797,
	-0.127737441217663,
	-0.126215877078991,
	-0.124694015942168,
	-0.123171861388281,
	-0.121649416999107,
	-0.120126686357102,
	-0.118603673045401,
	-0.117080380647801,
	-0.115556812748756,
	-0.114032972933368,
	-0.11250886478738,
	-0.110984491897164,
	-0.109459857849719,
	-0.107934966232654,
	-0.106409820634188,
	-0.104884424643136,
	-0.103358781848901,
	-0.101832895841467,
	-0.100306770211393,
	-0.0987804085498001,
	-0.0972538144483644,
	-0.0957269914993082,
	-0.094199943295394,
	-0.092672673429914,
	-0.0911451854966815,
	-0.0896174830900233,
	-0.0880895698047716,
	-0.0865614492362521,
	-0.085033124980281,
	-0.083504600633153,
	-0.0819758797916335,
	-0.0804469660529512,
	-0.0789178630147859,
	-0.0773885742752659,
	-0.0758591034329551,
	-0.0743294540868463,
	-0.072799629836352,
	-0.0712696342812975,
	-0.0697394710219082,
	-0.0682091436588071,
	-0.0666786557930022,
	-0.0651480110258793,
	-0.0636172129591943,
	-0.0620862651950611,
	-0.0605551713359486,
	-0.0590239349846686,
	-0.0574925597443681,
	-0.0559610492185209,
	-0.0544294070109202,
	-0.0528976367256662,
	-0.0513657419671634,
	-0.0498337263401079,
	-0.0483015934494806,
	-0.046769346900539,
	-0.0452369902988056,
	-0.0437045272500643,
	-0.0421719613603486,
	-0.0406392962359343,
	-0.0391065354833302,
	-0.0375736827092716,
	-0.0360407415207072,
	-0.0345077155247965,
	-0.0329746083288979,
	-0.0314414235405607,
	-0.0299081647675177,
	-0.0283748356176731,
	-0.0268414396990994,
	-0.0253079806200253,
	-0.0237744619888281,
	-0.0222408874140253,
	-0.020707260504267,
	-0.0191735848683235,
	-0.0176398641150828,
	-0.0161061018535379,
	-0.0145723016927795,
	-0.0130384672419885,
	-0.0115046021104237,
	-0.00997070990741888,
	-0.00843679424237049,
	-0.00690285872473028,
	-0.00536890696399671,
	-0.00383494256970732,
	-0.00230096915142674,
	-0.000766990318743474
  		 )
       );

  port (
    -- Sequential logic inside this unit
    iClk         : in std_ulogic;
    inResetAsync : in std_ulogic;

    -- Phase steps determining the frequency to be generated
    iPhaseIncrement : in natural range 0 to 2**(gPhaseResolution-1)-1;

    -- Sample rate sync strobe signal
    iSampleStrobe : in std_ulogic;

    -- Parallel digital audio data protocol
    oVal : out std_ulogic;
    oD   : out aAudioData(0 downto -(gAudioBitWidth-1)));

begin

  -- Assure that gWaveTable is of the form 2**n!
  assert 2**LogDualis(gWaveTable'length) = gWaveTable'length
    report "gWaveTable must have 2**n entries, but has " &
           natural'image(gWaveTable'length)
    severity error;
  
  -- Assure phase resolution is equal to or higher than the number of ROM address bits
  assert gPhaseResolution >= LogDualis(gWaveTable'length)
    report "gPhaseResolution is lower than the number of address bits necessary to address each table entry in gWaveTable"
    severity error;
  
  -- Assure that no more than the complete phase register is dithered
  assert gNrOfPhaseDitherBits <= gPhaseResolution
    report "Cannot dither more bits than those used to address the wave table"
    severity error;
  
  -- Warn if phase dithering is not set to the optimum (see comment for gNrOfPhaseDitherBits)
  assert gNrOfPhaseDitherBits = (gPhaseResolution - LogDualis(gWaveTable'length))
    report "Number of phase dithering bits deviates from ideal value " &
           "(is "       & integer'image(gNrOfPhaseDitherBits)                            & " bits," &
           " expected " & integer'image(gPhaseResolution - LogDualis(gWaveTable'length)) & " bits)"
    severity warning;
  
end DspDds;
