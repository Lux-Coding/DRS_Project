library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.Global.all;
use work.DefinitionsCodec.all;
use work.ParamCodec.all;
use work.DefinitionsFsk.all;
use work.InterfaceFunctions.all;

entity DataDetector is
    generic (
        gClkFrequency       : integer := cDefaultClkFrequency;
        gDistanceOne_us     : integer := 900;
        gDistanceTwo_us     : integer := 99900;
        gDistanceThree_us   : integer := 499900;
        gDistanceFour_us    : integer := 999900;
        gBaudRate           : integer := 9600;
        gDetectData         : std_ulogic_vector(7 downto 0) := x"0A";
        gDetectCycleLength  : integer := 4
    );
    port (
        iClk            :  in std_ulogic;
        inResetAsync    :  in std_ulogic;
        -- input data
        iData           :  in std_ulogic;
        iDistanceSelect :  in std_ulogic_vector(1 downto 0);
        -- data byte detected
        oByteDetected   : out std_ulogic;
        oSegDistance    : out std_logic_vector(6 downto 0)  -- active low
    );
end entity DataDetector;
