--------------------------------------------------------------------------------
-- Title       : Parameter definitions for FSK modem
-- Project     : FPGA Based Digital Signal Processing
--               FH O� Hagenberg/HSD, SCD5
--------------------------------------------------------------------------------
-- RevCtrl     : $Id: DefinitionsFsk-p.vhd 733 2017-12-04 02:28:35Z mroland $
-- Authors     : Michael Roland, Hagenberg/Austria, Copyright (c) 2015-2017
--------------------------------------------------------------------------------
-- Description : Channel frequency definitions and filter coefficients for FSK
--               modem
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.Global.all;

package DefinitionsFsk is

  type aTxFrequencySet is record
    Frequency0 : real;
    Frequency1 : real;
  end record;
  
  type aPhaseIncrementSet is record
    PhaseIncrement0 : natural;
    PhaseIncrement1 : natural;
  end record;
  
  type aSetOfTxChannels is array (natural range <>) of aTxFrequencySet;
  type aSetOfPhaseIncrements is array (natural range <>) of aPhaseIncrementSet;
  
  constant cFskFilterCoefWidth : natural := 16;
  constant cFskBandpassOrder   : natural := 257;
  constant cFskLowpassOrder    : natural := 74;

  constant cFskBandpassOrderDRS : natural := 190;
  constant cFskLowpassOrderDRS  : natural := 127;
  
  type aRxBandpassSet is record
    Bandpass0 : aSetOfFactors(0 to cFskBandpassOrderDRS);
    Bandpass1 : aSetOfFactors(0 to cFskBandpassOrderDRS);
  end record;

  type aSetOfRxBandpasses is array (natural range <>) of aRxBandpassSet;

  --constant cLowpass : aSetOfFactors(0 to cFskLowpassOrder) := (-0.000152587890625000, -9.15527343750000e-05, -9.15527343750000e-05, -9.15527343750000e-05, -6.10351562500000e-05, 0.0,  0.000122070312500000, 0.000274658203125000, 0.000488281250000000, 0.000793457031250000, 0.00119018554687500, 0.00167846679687500, 0.00231933593750000, 0.00305175781250000, 0.00396728515625000, 0.00503540039062500, 0.00622558593750000, 0.00762939453125000, 0.00915527343750000, 0.0108642578125000, 0.0127258300781250, 0.0147094726562500, 0.0168151855468750, 0.0190124511718750, 0.0212707519531250, 0.0235900878906250, 0.0258789062500000, 0.0281677246093750, 0.0303955078125000, 0.0325012207031250, 0.0344543457031250, 0.0362548828125000, 0.0378417968750000, 0.0391540527343750, 0.0402221679687500, 0.0410156250000000, 0.0414733886718750, 0.0416564941406250, 0.0414733886718750, 0.0410156250000000, 0.0402221679687500, 0.0391540527343750, 0.0378417968750000, 0.0362548828125000, 0.0344543457031250, 0.0325012207031250, 0.0303955078125000, 0.0281677246093750, 0.0258789062500000, 0.0235900878906250, 0.0212707519531250, 0.0190124511718750, 0.0168151855468750, 0.0147094726562500, 0.0127258300781250, 0.0108642578125000, 0.00915527343750000, 0.00762939453125000, 0.00622558593750000, 0.00503540039062500, 0.00396728515625000, 0.00305175781250000, 0.00231933593750000, 0.00167846679687500, 0.00119018554687500, 0.000793457031250000, 0.000488281250000000, 0.000274658203125000, 0.000122070312500000, 0.0,  -6.10351562500000e-05, -9.15527343750000e-05, -9.15527343750000e-05, -9.15527343750000e-05, -0.000152587890625000);

  constant cZeroBandpass : aSetOfFactors(0 to cFskBandpassOrderDRS) := (others => 0.0);

  constant cBandpass0Ch4 : aSetOfFactors(0 to cFskBandpassOrder) := (0.000916487968635350, 0.00203491092085189, -0.000590559011667039, -0.000354187586647468, -0.000780187537689414, -2.03384678617515e-05, 0.000694058720405891, 0.000853905489978949, 0.000118733222181907, -0.000823972325463847, -0.00103674827648814, -0.000201567343639594, 0.000941369069995207, 0.00124788970816623, 0.000304473701964881, -0.00105709684782540, -0.00148149243905214, -0.000431818748815704, 0.00116975748798141, 0.00173790182645744, 0.000586544983405864, -0.00127675427112592, -0.00201672839032318, -0.000771631063308161, 0.00137324726263239, 0.00231426508903349, 0.000986500332990503, -0.00145785299306605, -0.00263069603050938, -0.00123514602943768, 0.00152494191014539, 0.00296299501551174, 0.00151837806840317, -0.00157210842247685, -0.00330930181364335, -0.00183681883013199, 0.00159547427536924, 0.00366560070604853, 0.00219036347616303, -0.00159068330280919, -0.00402836976636600, -0.00258035771529688, 0.00155417184389778, 0.00439469978032757, 0.00300538472048231, -0.00148362010288037, -0.00475860148075850, -0.00346302886432834, 0.00137466322286556, 0.00511621276525590, 0.00395372370258572, -0.00122533632515662, -0.00546305439520559, -0.00447268407161426, 0.00103295647030899, 0.00579271535983805, 0.00501901976050332, -0.000795305471094868, -0.00610185740252455, -0.00558734745299377, 0.000511713802636828, 0.00638331078550669, 0.00617487562071629, -0.000180258367899253, -0.00663384555304851, -0.00677558336962589, -0.000198306322031002, 0.00684669503185135, 0.00738560264416012, 0.000623172049577571, -0.00701876036947186, -0.00799769536823997, -0.00109386241361189, 0.00714461879743551, 0.00860722996474740, 0.00160720865894132, -0.00722053377020737, -0.00920748328911600, -0.00216162878237644, 0.00724416571808825, 0.00979127659709388, 0.00275328021509339, -0.00721143862623890, -0.0103536348757699, -0.00337757909947203, 0.00712008658792456, 0.0108875109806534, 0.00403052892552971, -0.00696991697794312, -0.0113856176871422, -0.00470694939786154, 0.00675946123788833, 0.0118429190983579, 0.00540036136495933, -0.00648857055040806, -0.0122537439730605, -0.00610391105508545, 0.00615815390715540, 0.0126120726600280, 0.00681221560485166, -0.00577074671389308, -0.0129131238548969, -0.00751765918163146, 0.00532869940733876, 0.0131524549469569, 0.00821332485198605, -0.00483481486129901, -0.0133270350358977, -0.00889180232883397, 0.00429365094742298, 0.0134337071638497, 0.00954607497784231, -0.00370940869980489, -0.0134710196608538, -0.0101690738155750, 0.00308806286528727, 0.0134370361593299, 0.0107543748948239, -0.00243518488286462, -0.0133320027593651, -0.0112956641839960, 0.00175758958472457, 0.0131562444968423, 0.0117868094910609, -0.00106181370082753, -0.0129110880563249, -0.0122228997682831, 0.000355160256794235, 0.0125989169088260, 0.0125989169088260, 0.000355160256794235, -0.0122228997682831, -0.0129110880563249, -0.00106181370082753, 0.0117868094910609, 0.0131562444968423, 0.00175758958472457, -0.0112956641839960, -0.0133320027593651, -0.00243518488286462, 0.0107543748948239, 0.0134370361593299, 0.00308806286528727, -0.0101690738155750, -0.0134710196608538, -0.00370940869980489, 0.00954607497784231, 0.0134337071638497, 0.00429365094742298, -0.00889180232883397, -0.0133270350358977, -0.00483481486129901, 0.00821332485198605, 0.0131524549469569, 0.00532869940733876, -0.00751765918163146, -0.0129131238548969, -0.00577074671389308, 0.00681221560485166, 0.0126120726600280, 0.00615815390715540, -0.00610391105508545, -0.0122537439730605, -0.00648857055040806, 0.00540036136495933, 0.0118429190983579, 0.00675946123788833, -0.00470694939786154, -0.0113856176871422, -0.00696991697794312, 0.00403052892552971, 0.0108875109806534, 0.00712008658792456, -0.00337757909947203, -0.0103536348757699, -0.00721143862623890, 0.00275328021509339, 0.00979127659709388, 0.00724416571808825, -0.00216162878237644, -0.00920748328911600, -0.00722053377020737, 0.00160720865894132, 0.00860722996474740, 0.00714461879743551, -0.00109386241361189, -0.00799769536823997, -0.00701876036947186, 0.000623172049577571, 0.00738560264416012, 0.00684669503185135, -0.000198306322031002, -0.00677558336962589, -0.00663384555304851, -0.000180258367899253, 0.00617487562071629, 0.00638331078550669, 0.000511713802636828, -0.00558734745299377, -0.00610185740252455, -0.000795305471094868, 0.00501901976050332, 0.00579271535983805, 0.00103295647030899, -0.00447268407161426, -0.00546305439520559, -0.00122533632515662, 0.00395372370258572, 0.00511621276525590, 0.00137466322286556, -0.00346302886432834, -0.00475860148075850, -0.00148362010288037, 0.00300538472048231, 0.00439469978032757, 0.00155417184389778, -0.00258035771529688, -0.00402836976636600, -0.00159068330280919, 0.00219036347616303, 0.00366560070604853, 0.00159547427536924, -0.00183681883013199, -0.00330930181364335, -0.00157210842247685, 0.00151837806840317, 0.00296299501551174, 0.00152494191014539, -0.00123514602943768, -0.00263069603050938, -0.00145785299306605, 0.000986500332990503, 0.00231426508903349, 0.00137324726263239, -0.000771631063308161, -0.00201672839032318, -0.00127675427112592, 0.000586544983405864, 0.00173790182645744, 0.00116975748798141, -0.000431818748815704, -0.00148149243905214, -0.00105709684782540, 0.000304473701964881, 0.00124788970816623, 0.000941369069995207, -0.000201567343639594, -0.00103674827648814, -0.000823972325463847, 0.000118733222181907, 0.000853905489978949, 0.000694058720405891, -2.03384678617515e-05, -0.000780187537689414, -0.000354187586647468, -0.000590559011667039, 0.00203491092085189, 0.000916487968635350);
  constant cBandpass1Ch4 : aSetOfFactors(0 to cFskBandpassOrder) := (0.000984652195063242, 0.00182188651736983, -0.00116961973741390, -1.86771168986534e-05, 0.000615718610693588, 0.000143915284337272, -0.000883381268895002, 0.000170226912954838, 0.000924089867889370, -0.000470325143262863, -0.000899347112849682, 0.000810034175889535, 0.000755892863967181, -0.00113978069115514, -0.000489834311421356, 0.00141899717141631, 0.000105712461137516, -0.00160374142646866, 0.000377418019644007, 0.00165133795278037, -0.000922748620553012, -0.00152987244591735, 0.00148140257954482, 0.00121912651063238, -0.00199171823133018, -0.000719783349164338, 0.00238882284776716, 5.22174355458773e-05, -0.00260748494292771, 0.000738645987471043, 0.00259459657723147, -0.00159067744189936, -0.00231567292390517, 0.00241734543798856, 0.00175582851478124, -0.00313183544893376, -0.000932474228861696, 0.00363980363449256, -0.000105931439641748, -0.00386023042978427, 0.00128362482037627, 0.00372868073678962, -0.00249626036346685, -0.00321360953453676, 0.00362604855930261, 0.00231667675692028, -0.00454659515792367, -0.00108287681563732, 0.00514113603911372, -0.000405601723228253, -0.00531042115673260, 0.00202847494005081, 0.00499006476574315, -0.00364006468293778, -0.00415738421706104, 0.00507893607588331, 0.00284160197078172, -0.00618668418796999, -0.00112219859995927, 0.00682107154595127, -0.000871687929707449, -0.00687560275113219, 0.00297427138697957, 0.00629045754792885, -0.00498902684307777, -0.00506574426823123, 0.00671571216818182, 0.00326441530979638, -0.00796356809262721, -0.00101232312478285, 0.00857564275331623, -0.00151232550122033, -0.00844317903774439, 0.00408901569909103, 0.00752404862234650, -0.00647717498773257, -0.00584924875091293, 0.00843808919048361, 0.00352571549419292, -0.00975927307991600, -0.000728416832607551, 0.0102742000063684, -0.00230813765584706, -0.00988695211905504, 0.00531484059581778, 0.00858108981167503, -0.00800979436178187, -0.00642709342467240, 0.0101253382285931, 0.00358047950655756, -0.0114345308636865, -0.000272266096523669, 0.0117788394652025, -0.00321580113542137, -0.0110807827010075, 0.00656780602476586, 0.00936050928726403, -0.00947019196046453, -0.00673513915147317, 0.0116391756055820, 0.00341054436592971, -0.0128483518600714, 0.000333110316193327, 0.0129543901182152, -0.00416704216482718, -0.0119137765556958, 0.00774535003333818, 0.00978627346025206, -0.0107333773994850, -0.00673876362631901, 0.0128468876722250, 0.00302315538371185, -0.0138714144986096, 0.00103581003119030, 0.0136941190955383, -0.00507932174440091, -0.0123075117579959, 0.00874034667493386, 0.00981868315414162, -0.0116838829641630, -0.00643664625621716, 0.0136353948920964, 0.00245654792558669, -0.0144096444642028, 0.00176944199604945, 0.0139281859195889, -0.00586304040430037, -0.0122274991413658, 0.00945663775897771, 0.00945663775897771, -0.0122274991413658, -0.00586304040430037, 0.0139281859195889, 0.00176944199604945, -0.0144096444642028, 0.00245654792558669, 0.0136353948920964, -0.00643664625621716, -0.0116838829641630, 0.00981868315414162, 0.00874034667493386, -0.0123075117579959, -0.00507932174440091, 0.0136941190955383, 0.00103581003119030, -0.0138714144986096, 0.00302315538371185, 0.0128468876722250, -0.00673876362631901, -0.0107333773994850, 0.00978627346025206, 0.00774535003333818, -0.0119137765556958, -0.00416704216482718, 0.0129543901182152, 0.000333110316193327, -0.0128483518600714, 0.00341054436592971, 0.0116391756055820, -0.00673513915147317, -0.00947019196046453, 0.00936050928726403, 0.00656780602476586, -0.0110807827010075, -0.00321580113542137, 0.0117788394652025, -0.000272266096523669, -0.0114345308636865, 0.00358047950655756, 0.0101253382285931, -0.00642709342467240, -0.00800979436178187, 0.00858108981167503, 0.00531484059581778, -0.00988695211905504, -0.00230813765584706, 0.0102742000063684, -0.000728416832607551, -0.00975927307991600, 0.00352571549419292, 0.00843808919048361, -0.00584924875091293, -0.00647717498773257, 0.00752404862234650, 0.00408901569909103, -0.00844317903774439, -0.00151232550122033, 0.00857564275331623, -0.00101232312478285, -0.00796356809262721, 0.00326441530979638, 0.00671571216818182, -0.00506574426823123, -0.00498902684307777, 0.00629045754792885, 0.00297427138697957, -0.00687560275113219, -0.000871687929707449, 0.00682107154595127, -0.00112219859995927, -0.00618668418796999, 0.00284160197078172, 0.00507893607588331, -0.00415738421706104, -0.00364006468293778, 0.00499006476574315, 0.00202847494005081, -0.00531042115673260, -0.000405601723228253, 0.00514113603911372, -0.00108287681563732, -0.00454659515792367, 0.00231667675692028, 0.00362604855930261, -0.00321360953453676, -0.00249626036346685, 0.00372868073678962, 0.00128362482037627, -0.00386023042978427, -0.000105931439641748, 0.00363980363449256, -0.000932474228861696, -0.00313183544893376, 0.00175582851478124, 0.00241734543798856, -0.00231567292390517, -0.00159067744189936, 0.00259459657723147, 0.000738645987471043, -0.00260748494292771, 5.22174355458773e-05, 0.00238882284776716, -0.000719783349164338, -0.00199171823133018, 0.00121912651063238, 0.00148140257954482, -0.00152987244591735, -0.000922748620553012, 0.00165133795278037, 0.000377418019644007, -0.00160374142646866, 0.000105712461137516, 0.00141899717141631, -0.000489834311421356, -0.00113978069115514, 0.000755892863967181, 0.000810034175889535, -0.000899347112849682, -0.000470325143262863, 0.000924089867889370, 0.000170226912954838, -0.000883381268895002, 0.000143915284337272, 0.000615718610693588, -1.86771168986534e-05, -0.00116961973741390, 0.00182188651736983, 0.000984652195063242);

  constant cBandpass0Ch7 : aSetOfFactors(0 to cFskBandpassOrder) := (0.000896390789053966, 0.00200843767241717, -0.000673148718857462, -0.000433482166009556, -0.000618277023117879, 0.000327266688385479, 0.000847716575178528, 0.000462837843965778, -0.000565211830101954, -0.00102675869816148, -0.000298285532341100, 0.000885194955836250, 0.00113407437982955, 3.53870081485537e-05, -0.00123251844787957, -0.00114990481132625, 0.000332230857995906, 0.00157188259781267, 0.00104515716878642, -0.000794616157609980, -0.00186219600121912, -0.000795326032082708, 0.00132919082597881, 0.00205845788804461, 0.000386281866301376, -0.00190005288044732, -0.00211541363672818, 0.000179997611588692, 0.00245514393593316, 0.00198902456360711, -0.000887944290646646, -0.00293765400917211, -0.00165066418727747, 0.00170026893712578, 0.00328366111287915, 0.00108286857655443, -0.00256532585302284, -0.00343058822945577, -0.000287942534725186, 0.00341357021291263, 0.00332265767176740, -0.000707298090309838, -0.00416493464901705, -0.00292044477626431, 0.00185388358036924, 0.00473564189595204, 0.00220239649499888, -0.00308103707415937, -0.00504190216627546, -0.00117370294359889, 0.00429633683112024, 0.00501330210947055, -0.000129941937033568, -0.00539701785578929, -0.00459659204609373, 0.00164667808831575, 0.00627305263908726, 0.00376644494504611, -0.00328247561604150, -0.00682085557579762, -0.00252944791239369, 0.00492509283308027, 0.00694883929844901, 0.000927442560714108, -0.00644305035901050, -0.00659233637994627, 0.000961119722211973, 0.00770279835857169, 0.00571670455614960, -0.00302436476954302, -0.00857470581099482, -0.00432904739256239, 0.00512545418694585, 0.00894760986711145, 0.00247659973576025, -0.00710682741458246, -0.00874062965080589, -0.000251140962151990, 0.00880806346931790, 0.00790951565606855, -0.00221710137334233, -0.0100759406930370, -0.00645803638860809, 0.00476838131718411, 0.0107761642807665, 0.00443920024641677, -0.00722211997602278, -0.0108110897560823, -0.00195358104515732, 0.00939138142303362, 0.0101269197537192, -0.000854128987614965, -0.0110984147168175, -0.00872107657222194, 0.00380347359699762, 0.0121900372852488, 0.00664658139192184, -0.00669283953621046, -0.0125503132581594, -0.00401103385992828, 0.00931381525988918, 0.0121119326598343, 0.000971151384250557, -0.0114673891666252, -0.0108655276533346, 0.00227945522873917, 0.0129806626962516, 0.00886217543337185, -0.00552261039922913, -0.0137206791071698, -0.00621162627207788, 0.00853213991436139, 0.0136087570842718, 0.00307547036424719, -0.0110922242044333, -0.0126261307325182, 0.000343567135611963, 0.0130141768433426, 0.0108183136787658, -0.00381743229649020, -0.0141515178360400, -0.00829263965045894, 0.00710887753756899, 0.0144136592686750, 0.00521075622979819, -0.00999109378249707, -0.0137719762758637, -0.00177707155511109, 0.0122641395424944, 0.0122641395424944, -0.00177707155511109, -0.0137719762758637, -0.00999109378249707, 0.00521075622979819, 0.0144136592686750, 0.00710887753756899, -0.00829263965045894, -0.0141515178360400, -0.00381743229649020, 0.0108183136787658, 0.0130141768433426, 0.000343567135611963, -0.0126261307325182, -0.0110922242044333, 0.00307547036424719, 0.0136087570842718, 0.00853213991436139, -0.00621162627207788, -0.0137206791071698, -0.00552261039922913, 0.00886217543337185, 0.0129806626962516, 0.00227945522873917, -0.0108655276533346, -0.0114673891666252, 0.000971151384250557, 0.0121119326598343, 0.00931381525988918, -0.00401103385992828, -0.0125503132581594, -0.00669283953621046, 0.00664658139192184, 0.0121900372852488, 0.00380347359699762, -0.00872107657222194, -0.0110984147168175, -0.000854128987614965, 0.0101269197537192, 0.00939138142303362, -0.00195358104515732, -0.0108110897560823, -0.00722211997602278, 0.00443920024641677, 0.0107761642807665, 0.00476838131718411, -0.00645803638860809, -0.0100759406930370, -0.00221710137334233, 0.00790951565606855, 0.00880806346931790, -0.000251140962151990, -0.00874062965080589, -0.00710682741458246, 0.00247659973576025, 0.00894760986711145, 0.00512545418694585, -0.00432904739256239, -0.00857470581099482, -0.00302436476954302, 0.00571670455614960, 0.00770279835857169, 0.000961119722211973, -0.00659233637994627, -0.00644305035901050, 0.000927442560714108, 0.00694883929844901, 0.00492509283308027, -0.00252944791239369, -0.00682085557579762, -0.00328247561604150, 0.00376644494504611, 0.00627305263908726, 0.00164667808831575, -0.00459659204609373, -0.00539701785578929, -0.000129941937033568, 0.00501330210947055, 0.00429633683112024, -0.00117370294359889, -0.00504190216627546, -0.00308103707415937, 0.00220239649499888, 0.00473564189595204, 0.00185388358036924, -0.00292044477626431, -0.00416493464901705, -0.000707298090309838, 0.00332265767176740, 0.00341357021291263, -0.000287942534725186, -0.00343058822945577, -0.00256532585302284, 0.00108286857655443, 0.00328366111287915, 0.00170026893712578, -0.00165066418727747, -0.00293765400917211, -0.000887944290646646, 0.00198902456360711, 0.00245514393593316, 0.000179997611588692, -0.00211541363672818, -0.00190005288044732, 0.000386281866301376, 0.00205845788804461, 0.00132919082597881, -0.000795326032082708, -0.00186219600121912, -0.000794616157609980, 0.00104515716878642, 0.00157188259781267, 0.000332230857995906, -0.00114990481132625, -0.00123251844787957, 3.53870081485537e-05, 0.00113407437982955, 0.000885194955836250, -0.000298285532341100, -0.00102675869816148, -0.000565211830101954, 0.000462837843965778, 0.000847716575178528, 0.000327266688385479, -0.000618277023117879, -0.000433482166009556, -0.000673148718857462, 0.00200843767241717, 0.000896390789053966);
  constant cBandpass1Ch7 : aSetOfFactors(0 to cFskBandpassOrder) := (0.00100117732473863, 0.00176208667045678, -0.00120832133240698, 0.000151816197899113, 0.000629947630700073, -0.000202380031268052, -0.000746422372222872, 0.000674665968172095, 0.000473237443887142, -0.000996525435755381, -2.48252458895707e-05, 0.00113523831007643, -0.000556644113237243, -0.000982981609199433, 0.00112474585590995, 0.000517324224030808, -0.00151296002523003, 0.000200395855363677, 0.00156967720408900, -0.00102165332053276, -0.00120717565734864, 0.00173659239244129, 0.000440745997270173, -0.00212435114814704, 0.000596722732286446, 0.00201388023879622, -0.00167041880477174, -0.00134306323634697, 0.00249330454980393, 0.000194596639540985, -0.00279748222127933, 0.00120035042608349, 0.00241116065635449, -0.00251037359680961, -0.00133032702619410, 0.00336766805923078, -0.000266784910346012, -0.00347594073137290, 0.00203272038996709, 0.00269619895816910, -0.00352499071466614, -0.00110785447927983, 0.00431217780281501, -0.000982034376964320, -0.00409352836219096, 0.00309276696630070, 0.00279592296742675, -0.00467685024651900, -0.000622763806924845, 0.00525887026348853, -0.00196795166645810, -0.00457044179608640, 0.00435625427807876, 0.00264411792864291, -0.00590470491236510, 0.000160815449045033, 0.00612566309732953, -0.00321854282458913, -0.00482496578904227, 0.00577333140558033, 0.00218312781304657, -0.00712576666427816, 0.00125748134143546, 0.00682031180674637, -0.00469772119041124, -0.00478264920390960, 0.00726797375142785, 0.00137683972969849, -0.00824457469073602, 0.00265261162160296, 0.00725180271654261, -0.00634327851164303, -0.00438395153128187, 0.00874380156731617, 0.000217585270770542, -0.00915789444246696, 0.00430005343425031, 0.00734121469947271, -0.00806576383510887, -0.00359584204454775, 0.0100927234750213, -0.00127170210699368, -0.00976795996863082, 0.00612351830527804, 0.00702928570079834, -0.00975628544535738, -0.00241594269701258, 0.0112031757977727, -0.00303410956375447, -0.00999179825874419, 0.00802158096717398, 0.00628554404937970, -0.0112957430784510, -0.000877202462785951, 0.0119718492435364, -0.00498181661765587, -0.00977165762338354, 0.00987487500369071, 0.00511530017581035, -0.0125659468242864, 0.000953016402187499, 0.0123152913002679, -0.00700148113796453, -0.00908364116856772, 0.0115563369671025, 0.00356117616848363, -0.0134615903452964, 0.00297482817980839, 0.0121804695235505, -0.00896540739701128, -0.00794117128331272, 0.0129439275692464, 0.00170228500519282, -0.0139019558291224, 0.00506704531553043, 0.0115496241159383, -0.0107416731339092, -0.00639691061018507, 0.0139331766502136, -0.000353655251677575, -0.0138393876065110, 0.00709646013237785, 0.0104451178177321, -0.0122079295803750, -0.00453813380661617, 0.0144482671218076, -0.00247953137073832, -0.0132639793312354, 0.00892900788428495, 0.00892900788428495, -0.0132639793312354, -0.00247953137073832, 0.0144482671218076, -0.00453813380661617, -0.0122079295803750, 0.0104451178177321, 0.00709646013237785, -0.0138393876065110, -0.000353655251677575, 0.0139331766502136, -0.00639691061018507, -0.0107416731339092, 0.0115496241159383, 0.00506704531553043, -0.0139019558291224, 0.00170228500519282, 0.0129439275692464, -0.00794117128331272, -0.00896540739701128, 0.0121804695235505, 0.00297482817980839, -0.0134615903452964, 0.00356117616848363, 0.0115563369671025, -0.00908364116856772, -0.00700148113796453, 0.0123152913002679, 0.000953016402187499, -0.0125659468242864, 0.00511530017581035, 0.00987487500369071, -0.00977165762338354, -0.00498181661765587, 0.0119718492435364, -0.000877202462785951, -0.0112957430784510, 0.00628554404937970, 0.00802158096717398, -0.00999179825874419, -0.00303410956375447, 0.0112031757977727, -0.00241594269701258, -0.00975628544535738, 0.00702928570079834, 0.00612351830527804, -0.00976795996863082, -0.00127170210699368, 0.0100927234750213, -0.00359584204454775, -0.00806576383510887, 0.00734121469947271, 0.00430005343425031, -0.00915789444246696, 0.000217585270770542, 0.00874380156731617, -0.00438395153128187, -0.00634327851164303, 0.00725180271654261, 0.00265261162160296, -0.00824457469073602, 0.00137683972969849, 0.00726797375142785, -0.00478264920390960, -0.00469772119041124, 0.00682031180674637, 0.00125748134143546, -0.00712576666427816, 0.00218312781304657, 0.00577333140558033, -0.00482496578904227, -0.00321854282458913, 0.00612566309732953, 0.000160815449045033, -0.00590470491236510, 0.00264411792864291, 0.00435625427807876, -0.00457044179608640, -0.00196795166645810, 0.00525887026348853, -0.000622763806924845, -0.00467685024651900, 0.00279592296742675, 0.00309276696630070, -0.00409352836219096, -0.000982034376964320, 0.00431217780281501, -0.00110785447927983, -0.00352499071466614, 0.00269619895816910, 0.00203272038996709, -0.00347594073137290, -0.000266784910346012, 0.00336766805923078, -0.00133032702619410, -0.00251037359680961, 0.00241116065635449, 0.00120035042608349, -0.00279748222127933, 0.000194596639540985, 0.00249330454980393, -0.00134306323634697, -0.00167041880477174, 0.00201388023879622, 0.000596722732286446, -0.00212435114814704, 0.000440745997270173, 0.00173659239244129, -0.00120717565734864, -0.00102165332053276, 0.00156967720408900, 0.000200395855363677, -0.00151296002523003, 0.000517324224030808, 0.00112474585590995, -0.000982981609199433, -0.000556644113237243, 0.00113523831007643, -2.48252458895707e-05, -0.000996525435755381, 0.000473237443887142, 0.000674665968172095, -0.000746422372222872, -0.000202380031268052, 0.000629947630700073, 0.000151816197899113, -0.00120832133240698, 0.00176208667045678, 0.00100117732473863);
  
  constant cBandpass0DRS : aSetOfFactors(0 to cFskBandpassOrderDRS) := (0.000026702880859375, 0.000125885009765625, -0.00037384033203125, -0.000698089599609375, 0.001049041748046875, -0.0016326904296875, 0.001739501953125, -0.0012359619140625, 0.000003814697265625, 0.001720428466796875, -0.00342559814453125, 0.00446319580078125, -0.0042877197265625, 0.0027008056640625, -0.000003814697265625, -0.0030517578125, 0.00548553466796875, -0.0064544677734375, 0.00559234619140625, -0.00316619873046875, 0.000003814697265625, 0.002819061279296875, -0.004398345947265625, 0.004375457763671875, -0.003070831298828125, 0.0012969970703125, 0.0, -0.000209808349609375, -0.000640869140625, 0.00191497802734375, -0.002655029296875, 0.002079010009765625, 0.0, -0.003009796142578125, 0.005809783935546875, -0.007198333740234375, 0.00646209716796875, -0.003734588623046875, 0.0, 0.00334930419921875, -0.005115509033203125, 0.00485992431640625, -0.0030975341796875, 0.00104522705078125, 0.0, 0.000667572021484375, -0.002742767333984375, 0.005001068115234375, -0.005863189697265625, 0.004207611083984375, 0.0, -0.005523681640625, 0.01032257080078125, -0.012416839599609375, 0.010822296142578125, -0.006069183349609375, 0.0, 0.005008697509765625, -0.0071563720703125, 0.00608062744140625, -0.003047943115234375, 0.000316619873046875, 0.0, 0.00289154052734375, -0.007900238037109375, 0.012401580810546875, -0.013423919677734375, 0.009151458740234375, 0.0, -0.01125335693359375, 0.0205078125, -0.024097442626953125, 0.0204925537109375, -0.011157989501953125, 0.0, 0.00833892822265625, -0.010700225830078125, 0.007053375244140625, -0.000701904296875, -0.003147125244140625, 0.0, 0.0113525390625, -0.02748870849609375, 0.0411376953125, -0.04392242431640625, 0.0301513671875, 0.0, -0.039371490478515625, 0.07553863525390625, -0.09497833251953125, 0.088199615478515625, -0.053836822509765625, 0.0, 0.0578765869140625, -0.10204315185546875, 0.11852264404296875, -0.10204315185546875, 0.0578765869140625, 0.0, -0.053836822509765625, 0.088199615478515625, -0.09497833251953125, 0.07553863525390625, -0.039371490478515625, 0.0, 0.0301513671875, -0.04392242431640625, 0.0411376953125, -0.02748870849609375, 0.0113525390625, 0.0, -0.003147125244140625, -0.000701904296875, 0.007053375244140625, -0.010700225830078125, 0.00833892822265625, 0.0, -0.011157989501953125, 0.0204925537109375, -0.024097442626953125, 0.0205078125, -0.01125335693359375, 0.0, 0.009151458740234375, -0.013423919677734375, 0.012401580810546875, -0.007900238037109375, 0.00289154052734375, 0.0, 0.000316619873046875, -0.003047943115234375, 0.00608062744140625, -0.0071563720703125, 0.005008697509765625, 0.0, -0.006069183349609375, 0.010822296142578125, -0.012416839599609375, 0.01032257080078125, -0.005523681640625, 0.0, 0.004207611083984375, -0.005863189697265625, 0.005001068115234375, -0.002742767333984375, 0.000667572021484375, 0.0, 0.00104522705078125, -0.0030975341796875, 0.00485992431640625, -0.005115509033203125, 0.00334930419921875, 0.0, -0.003734588623046875, 0.00646209716796875, -0.007198333740234375, 0.005809783935546875, -0.003009796142578125, 0.0, 0.002079010009765625, -0.002655029296875, 0.00191497802734375, -0.000640869140625, -0.000209808349609375, 0.0, 0.0012969970703125, -0.003070831298828125, 0.004375457763671875, -0.004398345947265625, 0.002819061279296875, 0.000003814697265625, -0.00316619873046875, 0.00559234619140625, -0.0064544677734375, 0.00548553466796875, -0.0030517578125, -0.000003814697265625, 0.0027008056640625, -0.0042877197265625, 0.00446319580078125, -0.00342559814453125, 0.001720428466796875, 0.000003814697265625, -0.0012359619140625, 0.001739501953125, -0.0016326904296875, 0.001049041748046875, -0.000698089599609375, -0.00037384033203125, 0.000125885009765625, 0.000026702880859375);
  constant cBandpass1DRS : aSetOfFactors(0 to cFskBandpassOrderDRS) := (0.00005340576171875, 0.000011444091796875, 0.000400543212890625, 0.000911712646484375, -0.00115203857421875, -0.000576019287109375, 0.001956939697265625, 0.0000152587890625, -0.002902984619140625, 0.001323699951171875, 0.0032958984375, -0.003162384033203125, -0.00275421142578125, 0.004993438720703125, 0.001129150390625, -0.00611114501953125, 0.0012359619140625, 0.005970001220703125, -0.003589630126953125, -0.004474639892578125, 0.005035400390625, 0.00215911865234375, -0.004978179931640625, 0.0, 0.00347137451171875, -0.000988006591796875, -0.00128173828125, 0.00029754638671875, -0.000415802001953125, 0.001773834228515625, 0.000598907470703125, -0.0041656494140625, 0.001007080078125, 0.005565643310546875, -0.00373077392578125, -0.005092620849609375, 0.006206512451171875, 0.00286102294921875, -0.007080078125, 0.0, 0.00579071044921875, -0.001857757568359375, -0.002971649169921875, 0.001476287841796875, 0.000240325927734375, 0.0012359619140625, 0.00061798095703125, -0.0050048828125, 0.001323699951171875, 0.007778167724609375, -0.005481719970703125, -0.0078125, 0.00991058349609375, 0.00475311279296875, -0.012256622314453125, 0.0, 0.011089324951171875, -0.0038299560546875, -0.006866455078125, 0.004299163818359375, 0.001953125, -0.000579833984375, 0.00048828125, -0.005786895751953125, 0.001781463623046875, 0.0114593505859375, -0.00861358642578125, -0.012943267822265625, 0.017192840576171875, 0.00861358642578125, -0.023227691650390625, 0.0, 0.0232086181640625, -0.00853729248046875, -0.01662445068359375, 0.011791229248046875, 0.006862640380859375, -0.006511688232421875, -0.000156402587890625, -0.0063018798828125, 0.002765655517578125, 0.020977020263671875, -0.01763916015625, -0.02909088134765625, 0.042171478271484375, 0.02307891845703125, -0.06836700439453125, 0.0, 0.085544586181640625, -0.036346435546875, -0.084674835205078125, 0.07613372802734375, 0.062412261962890625, -0.106937408447265625, -0.02298736572265625, 0.118518829345703125, -0.02298736572265625, -0.106937408447265625, 0.062412261962890625, 0.07613372802734375, -0.084674835205078125, -0.036346435546875, 0.085544586181640625, 0.0, -0.06836700439453125, 0.02307891845703125, 0.042171478271484375, -0.02909088134765625, -0.01763916015625, 0.020977020263671875, 0.002765655517578125, -0.0063018798828125, -0.000156402587890625, -0.006511688232421875, 0.006862640380859375, 0.011791229248046875, -0.01662445068359375, -0.00853729248046875, 0.0232086181640625, 0.0, -0.023227691650390625, 0.00861358642578125, 0.017192840576171875, -0.012943267822265625, -0.00861358642578125, 0.0114593505859375, 0.001781463623046875, -0.005786895751953125, 0.00048828125, -0.000579833984375, 0.001953125, 0.004299163818359375, -0.006866455078125, -0.0038299560546875, 0.011089324951171875, 0.0, -0.012256622314453125, 0.00475311279296875, 0.00991058349609375, -0.0078125, -0.005481719970703125, 0.007778167724609375, 0.001323699951171875, -0.0050048828125, 0.00061798095703125, 0.0012359619140625, 0.000240325927734375, 0.001476287841796875, -0.002971649169921875, -0.001857757568359375, 0.00579071044921875, 0.0, -0.007080078125, 0.00286102294921875, 0.006206512451171875, -0.005092620849609375, -0.00373077392578125, 0.005565643310546875, 0.001007080078125, -0.0041656494140625, 0.000598907470703125, 0.001773834228515625, -0.000415802001953125, 0.00029754638671875, -0.00128173828125, -0.000988006591796875, 0.00347137451171875, 0.0, -0.004978179931640625, 0.00215911865234375, 0.005035400390625, -0.004474639892578125, -0.003589630126953125, 0.005970001220703125, 0.0012359619140625, -0.00611114501953125, 0.001129150390625, 0.004993438720703125, -0.00275421142578125, -0.003162384033203125, 0.0032958984375, 0.001323699951171875, -0.002902984619140625, 0.0000152587890625, 0.001956939697265625, -0.000576019287109375, -0.00115203857421875, 0.000911712646484375, 0.000400543212890625, 0.000011444091796875, 0.00005340576171875);
  constant cLowpassDRS   : aSetOfFactors(0 to cFskLowpassOrderDRS) := (-0.0009632110595703125, -0.00006103515625, -0.00005245208740234375, -0.00003528594970703125, -0.00001049041748046875, 0.00002384185791015625, 0.00006866455078125, 0.00012493133544921875, 0.0001926422119140625, 0.0002727508544921875, 0.00036716461181640625, 0.00047588348388671875, 0.0006008148193359375, 0.0007419586181640625, 0.0009002685546875, 0.0010776519775390625, 0.00127410888671875, 0.0014896392822265625, 0.0017242431640625, 0.00198268890380859375, 0.0022602081298828125, 0.002559661865234375, 0.00288105010986328125, 0.00322437286376953125, 0.003589630126953125, 0.0039768218994140625, 0.0043849945068359375, 0.00481510162353515625, 0.0052642822265625, 0.005733489990234375, 0.006221771240234375, 0.00672817230224609375, 0.0072498321533203125, 0.0077877044677734375, 0.00833797454833984375, 0.00890064239501953125, 0.0094738006591796875, 0.0100555419921875, 0.01064395904541015625, 0.01123523712158203125, 0.01183032989501953125, 0.012424468994140625, 0.0130157470703125, 0.01360225677490234375, 0.01418209075927734375, 0.01475238800048828125, 0.01530933380126953125, 0.01585292816162109375, 0.0163784027099609375, 0.01688480377197265625, 0.01736927032470703125, 0.01782989501953125, 0.0182647705078125, 0.0186710357666015625, 0.019046783447265625, 0.019390106201171875, 0.01970005035400390625, 0.01997470855712890625, 0.02021312713623046875, 0.02041339874267578125, 0.0205745697021484375, 0.0206966400146484375, 0.02077770233154296875, 0.0208187103271484375, 0.0208187103271484375, 0.02077770233154296875, 0.0206966400146484375, 0.0205745697021484375, 0.02041339874267578125, 0.02021312713623046875, 0.01997470855712890625, 0.01970005035400390625, 0.019390106201171875, 0.019046783447265625, 0.0186710357666015625, 0.0182647705078125, 0.01782989501953125, 0.01736927032470703125, 0.01688480377197265625, 0.0163784027099609375, 0.01585292816162109375, 0.01530933380126953125, 0.01475238800048828125, 0.01418209075927734375, 0.01360225677490234375, 0.0130157470703125, 0.012424468994140625, 0.01183032989501953125, 0.01123523712158203125, 0.01064395904541015625, 0.0100555419921875, 0.0094738006591796875, 0.00890064239501953125, 0.00833797454833984375, 0.0077877044677734375, 0.0072498321533203125, 0.00672817230224609375, 0.006221771240234375, 0.005733489990234375, 0.0052642822265625, 0.00481510162353515625, 0.0043849945068359375, 0.0039768218994140625, 0.003589630126953125, 0.00322437286376953125, 0.00288105010986328125, 0.002559661865234375, 0.0022602081298828125, 0.00198268890380859375, 0.0017242431640625, 0.0014896392822265625, 0.00127410888671875, 0.0010776519775390625, 0.0009002685546875, 0.0007419586181640625, 0.0006008148193359375, 0.00047588348388671875, 0.00036716461181640625, 0.0002727508544921875, 0.0001926422119140625, 0.00012493133544921875, 0.00006866455078125, 0.00002384185791015625, -0.00001049041748046875, -0.00003528594970703125, -0.00005245208740234375, -0.00006103515625, -0.0009632110595703125);



end package DefinitionsFsk;


package body DefinitionsFsk is

  
end package body;
