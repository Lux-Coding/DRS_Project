-- Computer_System.vhd

-- Generated using ACDS version 16.0 211

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Computer_System is
	port (
		f2h_bootflags_boot_from_fpga_ready      : in    std_logic                     := '0';             -- f2h_bootflags.boot_from_fpga_ready
		f2h_bootflags_boot_from_fpga_on_failure : in    std_logic                     := '0';             --              .boot_from_fpga_on_failure
		fpga_reset_reset_n                      : out   std_logic;                                        --    fpga_reset.reset_n
		h2f_loan_io_in                          : out   std_logic_vector(66 downto 0);                    --   h2f_loan_io.in
		h2f_loan_io_out                         : in    std_logic_vector(66 downto 0) := (others => '0'); --              .out
		h2f_loan_io_oe                          : in    std_logic_vector(66 downto 0) := (others => '0'); --              .oe
		hps_io_hps_io_emac1_inst_TX_CLK         : out   std_logic;                                        --        hps_io.hps_io_emac1_inst_TX_CLK
		hps_io_hps_io_emac1_inst_TXD0           : out   std_logic;                                        --              .hps_io_emac1_inst_TXD0
		hps_io_hps_io_emac1_inst_TXD1           : out   std_logic;                                        --              .hps_io_emac1_inst_TXD1
		hps_io_hps_io_emac1_inst_TXD2           : out   std_logic;                                        --              .hps_io_emac1_inst_TXD2
		hps_io_hps_io_emac1_inst_TXD3           : out   std_logic;                                        --              .hps_io_emac1_inst_TXD3
		hps_io_hps_io_emac1_inst_RXD0           : in    std_logic                     := '0';             --              .hps_io_emac1_inst_RXD0
		hps_io_hps_io_emac1_inst_MDIO           : inout std_logic                     := '0';             --              .hps_io_emac1_inst_MDIO
		hps_io_hps_io_emac1_inst_MDC            : out   std_logic;                                        --              .hps_io_emac1_inst_MDC
		hps_io_hps_io_emac1_inst_RX_CTL         : in    std_logic                     := '0';             --              .hps_io_emac1_inst_RX_CTL
		hps_io_hps_io_emac1_inst_TX_CTL         : out   std_logic;                                        --              .hps_io_emac1_inst_TX_CTL
		hps_io_hps_io_emac1_inst_RX_CLK         : in    std_logic                     := '0';             --              .hps_io_emac1_inst_RX_CLK
		hps_io_hps_io_emac1_inst_RXD1           : in    std_logic                     := '0';             --              .hps_io_emac1_inst_RXD1
		hps_io_hps_io_emac1_inst_RXD2           : in    std_logic                     := '0';             --              .hps_io_emac1_inst_RXD2
		hps_io_hps_io_emac1_inst_RXD3           : in    std_logic                     := '0';             --              .hps_io_emac1_inst_RXD3
		hps_io_hps_io_qspi_inst_IO0             : inout std_logic                     := '0';             --              .hps_io_qspi_inst_IO0
		hps_io_hps_io_qspi_inst_IO1             : inout std_logic                     := '0';             --              .hps_io_qspi_inst_IO1
		hps_io_hps_io_qspi_inst_IO2             : inout std_logic                     := '0';             --              .hps_io_qspi_inst_IO2
		hps_io_hps_io_qspi_inst_IO3             : inout std_logic                     := '0';             --              .hps_io_qspi_inst_IO3
		hps_io_hps_io_qspi_inst_SS0             : out   std_logic;                                        --              .hps_io_qspi_inst_SS0
		hps_io_hps_io_qspi_inst_CLK             : out   std_logic;                                        --              .hps_io_qspi_inst_CLK
		hps_io_hps_io_sdio_inst_CMD             : inout std_logic                     := '0';             --              .hps_io_sdio_inst_CMD
		hps_io_hps_io_sdio_inst_D0              : inout std_logic                     := '0';             --              .hps_io_sdio_inst_D0
		hps_io_hps_io_sdio_inst_D1              : inout std_logic                     := '0';             --              .hps_io_sdio_inst_D1
		hps_io_hps_io_sdio_inst_CLK             : out   std_logic;                                        --              .hps_io_sdio_inst_CLK
		hps_io_hps_io_sdio_inst_D2              : inout std_logic                     := '0';             --              .hps_io_sdio_inst_D2
		hps_io_hps_io_sdio_inst_D3              : inout std_logic                     := '0';             --              .hps_io_sdio_inst_D3
		hps_io_hps_io_usb1_inst_D0              : inout std_logic                     := '0';             --              .hps_io_usb1_inst_D0
		hps_io_hps_io_usb1_inst_D1              : inout std_logic                     := '0';             --              .hps_io_usb1_inst_D1
		hps_io_hps_io_usb1_inst_D2              : inout std_logic                     := '0';             --              .hps_io_usb1_inst_D2
		hps_io_hps_io_usb1_inst_D3              : inout std_logic                     := '0';             --              .hps_io_usb1_inst_D3
		hps_io_hps_io_usb1_inst_D4              : inout std_logic                     := '0';             --              .hps_io_usb1_inst_D4
		hps_io_hps_io_usb1_inst_D5              : inout std_logic                     := '0';             --              .hps_io_usb1_inst_D5
		hps_io_hps_io_usb1_inst_D6              : inout std_logic                     := '0';             --              .hps_io_usb1_inst_D6
		hps_io_hps_io_usb1_inst_D7              : inout std_logic                     := '0';             --              .hps_io_usb1_inst_D7
		hps_io_hps_io_usb1_inst_CLK             : in    std_logic                     := '0';             --              .hps_io_usb1_inst_CLK
		hps_io_hps_io_usb1_inst_STP             : out   std_logic;                                        --              .hps_io_usb1_inst_STP
		hps_io_hps_io_usb1_inst_DIR             : in    std_logic                     := '0';             --              .hps_io_usb1_inst_DIR
		hps_io_hps_io_usb1_inst_NXT             : in    std_logic                     := '0';             --              .hps_io_usb1_inst_NXT
		hps_io_hps_io_spim1_inst_CLK            : out   std_logic;                                        --              .hps_io_spim1_inst_CLK
		hps_io_hps_io_spim1_inst_MOSI           : out   std_logic;                                        --              .hps_io_spim1_inst_MOSI
		hps_io_hps_io_spim1_inst_MISO           : in    std_logic                     := '0';             --              .hps_io_spim1_inst_MISO
		hps_io_hps_io_spim1_inst_SS0            : out   std_logic;                                        --              .hps_io_spim1_inst_SS0
		hps_io_hps_io_i2c0_inst_SDA             : inout std_logic                     := '0';             --              .hps_io_i2c0_inst_SDA
		hps_io_hps_io_i2c0_inst_SCL             : inout std_logic                     := '0';             --              .hps_io_i2c0_inst_SCL
		hps_io_hps_io_i2c1_inst_SDA             : inout std_logic                     := '0';             --              .hps_io_i2c1_inst_SDA
		hps_io_hps_io_i2c1_inst_SCL             : inout std_logic                     := '0';             --              .hps_io_i2c1_inst_SCL
		hps_io_hps_io_gpio_inst_GPIO09          : inout std_logic                     := '0';             --              .hps_io_gpio_inst_GPIO09
		hps_io_hps_io_gpio_inst_GPIO35          : inout std_logic                     := '0';             --              .hps_io_gpio_inst_GPIO35
		hps_io_hps_io_gpio_inst_GPIO40          : inout std_logic                     := '0';             --              .hps_io_gpio_inst_GPIO40
		hps_io_hps_io_gpio_inst_GPIO48          : inout std_logic                     := '0';             --              .hps_io_gpio_inst_GPIO48
		hps_io_hps_io_gpio_inst_GPIO61          : inout std_logic                     := '0';             --              .hps_io_gpio_inst_GPIO61
		hps_io_hps_io_gpio_inst_LOANIO49        : inout std_logic                     := '0';             --              .hps_io_gpio_inst_LOANIO49
		hps_io_hps_io_gpio_inst_LOANIO50        : inout std_logic                     := '0';             --              .hps_io_gpio_inst_LOANIO50
		hps_io_hps_io_gpio_inst_LOANIO53        : inout std_logic                     := '0';             --              .hps_io_gpio_inst_LOANIO53
		hps_io_hps_io_gpio_inst_LOANIO54        : inout std_logic                     := '0';             --              .hps_io_gpio_inst_LOANIO54
		hps_uart0_cts                           : in    std_logic                     := '0';             --     hps_uart0.cts
		hps_uart0_dsr                           : in    std_logic                     := '0';             --              .dsr
		hps_uart0_dcd                           : in    std_logic                     := '0';             --              .dcd
		hps_uart0_ri                            : in    std_logic                     := '0';             --              .ri
		hps_uart0_dtr                           : out   std_logic;                                        --              .dtr
		hps_uart0_rts                           : out   std_logic;                                        --              .rts
		hps_uart0_out1_n                        : out   std_logic;                                        --              .out1_n
		hps_uart0_out2_n                        : out   std_logic;                                        --              .out2_n
		hps_uart0_rxd                           : in    std_logic                     := '0';             --              .rxd
		hps_uart0_txd                           : out   std_logic;                                        --              .txd
		memory_mem_a                            : out   std_logic_vector(14 downto 0);                    --        memory.mem_a
		memory_mem_ba                           : out   std_logic_vector(2 downto 0);                     --              .mem_ba
		memory_mem_ck                           : out   std_logic;                                        --              .mem_ck
		memory_mem_ck_n                         : out   std_logic;                                        --              .mem_ck_n
		memory_mem_cke                          : out   std_logic;                                        --              .mem_cke
		memory_mem_cs_n                         : out   std_logic;                                        --              .mem_cs_n
		memory_mem_ras_n                        : out   std_logic;                                        --              .mem_ras_n
		memory_mem_cas_n                        : out   std_logic;                                        --              .mem_cas_n
		memory_mem_we_n                         : out   std_logic;                                        --              .mem_we_n
		memory_mem_reset_n                      : out   std_logic;                                        --              .mem_reset_n
		memory_mem_dq                           : inout std_logic_vector(31 downto 0) := (others => '0'); --              .mem_dq
		memory_mem_dqs                          : inout std_logic_vector(3 downto 0)  := (others => '0'); --              .mem_dqs
		memory_mem_dqs_n                        : inout std_logic_vector(3 downto 0)  := (others => '0'); --              .mem_dqs_n
		memory_mem_odt                          : out   std_logic;                                        --              .mem_odt
		memory_mem_dm                           : out   std_logic_vector(3 downto 0);                     --              .mem_dm
		memory_oct_rzqin                        : in    std_logic                     := '0';             --              .oct_rzqin
		system_clk_clk                          : in    std_logic                     := '0';             --    system_clk.clk
		system_reset_reset                      : in    std_logic                     := '0'              --  system_reset.reset
	);
end entity Computer_System;

architecture rtl of Computer_System is
	component Computer_System_ARM_A9_HPS is
		generic (
			F2S_Width : integer := 2;
			S2F_Width : integer := 2
		);
		port (
			h2f_loan_in                   : out   std_logic_vector(66 downto 0);                    -- in
			h2f_loan_out                  : in    std_logic_vector(66 downto 0) := (others => 'X'); -- out
			h2f_loan_oe                   : in    std_logic_vector(66 downto 0) := (others => 'X'); -- oe
			f2h_boot_from_fpga_ready      : in    std_logic                     := 'X';             -- boot_from_fpga_ready
			f2h_boot_from_fpga_on_failure : in    std_logic                     := 'X';             -- boot_from_fpga_on_failure
			uart0_cts                     : in    std_logic                     := 'X';             -- cts
			uart0_dsr                     : in    std_logic                     := 'X';             -- dsr
			uart0_dcd                     : in    std_logic                     := 'X';             -- dcd
			uart0_ri                      : in    std_logic                     := 'X';             -- ri
			uart0_dtr                     : out   std_logic;                                        -- dtr
			uart0_rts                     : out   std_logic;                                        -- rts
			uart0_out1_n                  : out   std_logic;                                        -- out1_n
			uart0_out2_n                  : out   std_logic;                                        -- out2_n
			uart0_rxd                     : in    std_logic                     := 'X';             -- rxd
			uart0_txd                     : out   std_logic;                                        -- txd
			mem_a                         : out   std_logic_vector(14 downto 0);                    -- mem_a
			mem_ba                        : out   std_logic_vector(2 downto 0);                     -- mem_ba
			mem_ck                        : out   std_logic;                                        -- mem_ck
			mem_ck_n                      : out   std_logic;                                        -- mem_ck_n
			mem_cke                       : out   std_logic;                                        -- mem_cke
			mem_cs_n                      : out   std_logic;                                        -- mem_cs_n
			mem_ras_n                     : out   std_logic;                                        -- mem_ras_n
			mem_cas_n                     : out   std_logic;                                        -- mem_cas_n
			mem_we_n                      : out   std_logic;                                        -- mem_we_n
			mem_reset_n                   : out   std_logic;                                        -- mem_reset_n
			mem_dq                        : inout std_logic_vector(31 downto 0) := (others => 'X'); -- mem_dq
			mem_dqs                       : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs
			mem_dqs_n                     : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs_n
			mem_odt                       : out   std_logic;                                        -- mem_odt
			mem_dm                        : out   std_logic_vector(3 downto 0);                     -- mem_dm
			oct_rzqin                     : in    std_logic                     := 'X';             -- oct_rzqin
			hps_io_emac1_inst_TX_CLK      : out   std_logic;                                        -- hps_io_emac1_inst_TX_CLK
			hps_io_emac1_inst_TXD0        : out   std_logic;                                        -- hps_io_emac1_inst_TXD0
			hps_io_emac1_inst_TXD1        : out   std_logic;                                        -- hps_io_emac1_inst_TXD1
			hps_io_emac1_inst_TXD2        : out   std_logic;                                        -- hps_io_emac1_inst_TXD2
			hps_io_emac1_inst_TXD3        : out   std_logic;                                        -- hps_io_emac1_inst_TXD3
			hps_io_emac1_inst_RXD0        : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD0
			hps_io_emac1_inst_MDIO        : inout std_logic                     := 'X';             -- hps_io_emac1_inst_MDIO
			hps_io_emac1_inst_MDC         : out   std_logic;                                        -- hps_io_emac1_inst_MDC
			hps_io_emac1_inst_RX_CTL      : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RX_CTL
			hps_io_emac1_inst_TX_CTL      : out   std_logic;                                        -- hps_io_emac1_inst_TX_CTL
			hps_io_emac1_inst_RX_CLK      : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RX_CLK
			hps_io_emac1_inst_RXD1        : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD1
			hps_io_emac1_inst_RXD2        : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD2
			hps_io_emac1_inst_RXD3        : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD3
			hps_io_qspi_inst_IO0          : inout std_logic                     := 'X';             -- hps_io_qspi_inst_IO0
			hps_io_qspi_inst_IO1          : inout std_logic                     := 'X';             -- hps_io_qspi_inst_IO1
			hps_io_qspi_inst_IO2          : inout std_logic                     := 'X';             -- hps_io_qspi_inst_IO2
			hps_io_qspi_inst_IO3          : inout std_logic                     := 'X';             -- hps_io_qspi_inst_IO3
			hps_io_qspi_inst_SS0          : out   std_logic;                                        -- hps_io_qspi_inst_SS0
			hps_io_qspi_inst_CLK          : out   std_logic;                                        -- hps_io_qspi_inst_CLK
			hps_io_sdio_inst_CMD          : inout std_logic                     := 'X';             -- hps_io_sdio_inst_CMD
			hps_io_sdio_inst_D0           : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D0
			hps_io_sdio_inst_D1           : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D1
			hps_io_sdio_inst_CLK          : out   std_logic;                                        -- hps_io_sdio_inst_CLK
			hps_io_sdio_inst_D2           : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D2
			hps_io_sdio_inst_D3           : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D3
			hps_io_usb1_inst_D0           : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D0
			hps_io_usb1_inst_D1           : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D1
			hps_io_usb1_inst_D2           : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D2
			hps_io_usb1_inst_D3           : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D3
			hps_io_usb1_inst_D4           : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D4
			hps_io_usb1_inst_D5           : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D5
			hps_io_usb1_inst_D6           : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D6
			hps_io_usb1_inst_D7           : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D7
			hps_io_usb1_inst_CLK          : in    std_logic                     := 'X';             -- hps_io_usb1_inst_CLK
			hps_io_usb1_inst_STP          : out   std_logic;                                        -- hps_io_usb1_inst_STP
			hps_io_usb1_inst_DIR          : in    std_logic                     := 'X';             -- hps_io_usb1_inst_DIR
			hps_io_usb1_inst_NXT          : in    std_logic                     := 'X';             -- hps_io_usb1_inst_NXT
			hps_io_spim1_inst_CLK         : out   std_logic;                                        -- hps_io_spim1_inst_CLK
			hps_io_spim1_inst_MOSI        : out   std_logic;                                        -- hps_io_spim1_inst_MOSI
			hps_io_spim1_inst_MISO        : in    std_logic                     := 'X';             -- hps_io_spim1_inst_MISO
			hps_io_spim1_inst_SS0         : out   std_logic;                                        -- hps_io_spim1_inst_SS0
			hps_io_i2c0_inst_SDA          : inout std_logic                     := 'X';             -- hps_io_i2c0_inst_SDA
			hps_io_i2c0_inst_SCL          : inout std_logic                     := 'X';             -- hps_io_i2c0_inst_SCL
			hps_io_i2c1_inst_SDA          : inout std_logic                     := 'X';             -- hps_io_i2c1_inst_SDA
			hps_io_i2c1_inst_SCL          : inout std_logic                     := 'X';             -- hps_io_i2c1_inst_SCL
			hps_io_gpio_inst_GPIO09       : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO09
			hps_io_gpio_inst_GPIO35       : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO35
			hps_io_gpio_inst_GPIO40       : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO40
			hps_io_gpio_inst_GPIO48       : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO48
			hps_io_gpio_inst_GPIO61       : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO61
			hps_io_gpio_inst_LOANIO49     : inout std_logic                     := 'X';             -- hps_io_gpio_inst_LOANIO49
			hps_io_gpio_inst_LOANIO50     : inout std_logic                     := 'X';             -- hps_io_gpio_inst_LOANIO50
			hps_io_gpio_inst_LOANIO53     : inout std_logic                     := 'X';             -- hps_io_gpio_inst_LOANIO53
			hps_io_gpio_inst_LOANIO54     : inout std_logic                     := 'X';             -- hps_io_gpio_inst_LOANIO54
			h2f_rst_n                     : out   std_logic;                                        -- reset_n
			h2f_axi_clk                   : in    std_logic                     := 'X';             -- clk
			h2f_AWID                      : out   std_logic_vector(11 downto 0);                    -- awid
			h2f_AWADDR                    : out   std_logic_vector(29 downto 0);                    -- awaddr
			h2f_AWLEN                     : out   std_logic_vector(3 downto 0);                     -- awlen
			h2f_AWSIZE                    : out   std_logic_vector(2 downto 0);                     -- awsize
			h2f_AWBURST                   : out   std_logic_vector(1 downto 0);                     -- awburst
			h2f_AWLOCK                    : out   std_logic_vector(1 downto 0);                     -- awlock
			h2f_AWCACHE                   : out   std_logic_vector(3 downto 0);                     -- awcache
			h2f_AWPROT                    : out   std_logic_vector(2 downto 0);                     -- awprot
			h2f_AWVALID                   : out   std_logic;                                        -- awvalid
			h2f_AWREADY                   : in    std_logic                     := 'X';             -- awready
			h2f_WID                       : out   std_logic_vector(11 downto 0);                    -- wid
			h2f_WDATA                     : out   std_logic_vector(63 downto 0);                    -- wdata
			h2f_WSTRB                     : out   std_logic_vector(7 downto 0);                     -- wstrb
			h2f_WLAST                     : out   std_logic;                                        -- wlast
			h2f_WVALID                    : out   std_logic;                                        -- wvalid
			h2f_WREADY                    : in    std_logic                     := 'X';             -- wready
			h2f_BID                       : in    std_logic_vector(11 downto 0) := (others => 'X'); -- bid
			h2f_BRESP                     : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- bresp
			h2f_BVALID                    : in    std_logic                     := 'X';             -- bvalid
			h2f_BREADY                    : out   std_logic;                                        -- bready
			h2f_ARID                      : out   std_logic_vector(11 downto 0);                    -- arid
			h2f_ARADDR                    : out   std_logic_vector(29 downto 0);                    -- araddr
			h2f_ARLEN                     : out   std_logic_vector(3 downto 0);                     -- arlen
			h2f_ARSIZE                    : out   std_logic_vector(2 downto 0);                     -- arsize
			h2f_ARBURST                   : out   std_logic_vector(1 downto 0);                     -- arburst
			h2f_ARLOCK                    : out   std_logic_vector(1 downto 0);                     -- arlock
			h2f_ARCACHE                   : out   std_logic_vector(3 downto 0);                     -- arcache
			h2f_ARPROT                    : out   std_logic_vector(2 downto 0);                     -- arprot
			h2f_ARVALID                   : out   std_logic;                                        -- arvalid
			h2f_ARREADY                   : in    std_logic                     := 'X';             -- arready
			h2f_RID                       : in    std_logic_vector(11 downto 0) := (others => 'X'); -- rid
			h2f_RDATA                     : in    std_logic_vector(63 downto 0) := (others => 'X'); -- rdata
			h2f_RRESP                     : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- rresp
			h2f_RLAST                     : in    std_logic                     := 'X';             -- rlast
			h2f_RVALID                    : in    std_logic                     := 'X';             -- rvalid
			h2f_RREADY                    : out   std_logic;                                        -- rready
			f2h_axi_clk                   : in    std_logic                     := 'X';             -- clk
			f2h_AWID                      : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- awid
			f2h_AWADDR                    : in    std_logic_vector(31 downto 0) := (others => 'X'); -- awaddr
			f2h_AWLEN                     : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- awlen
			f2h_AWSIZE                    : in    std_logic_vector(2 downto 0)  := (others => 'X'); -- awsize
			f2h_AWBURST                   : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- awburst
			f2h_AWLOCK                    : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- awlock
			f2h_AWCACHE                   : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- awcache
			f2h_AWPROT                    : in    std_logic_vector(2 downto 0)  := (others => 'X'); -- awprot
			f2h_AWVALID                   : in    std_logic                     := 'X';             -- awvalid
			f2h_AWREADY                   : out   std_logic;                                        -- awready
			f2h_AWUSER                    : in    std_logic_vector(4 downto 0)  := (others => 'X'); -- awuser
			f2h_WID                       : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- wid
			f2h_WDATA                     : in    std_logic_vector(63 downto 0) := (others => 'X'); -- wdata
			f2h_WSTRB                     : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- wstrb
			f2h_WLAST                     : in    std_logic                     := 'X';             -- wlast
			f2h_WVALID                    : in    std_logic                     := 'X';             -- wvalid
			f2h_WREADY                    : out   std_logic;                                        -- wready
			f2h_BID                       : out   std_logic_vector(7 downto 0);                     -- bid
			f2h_BRESP                     : out   std_logic_vector(1 downto 0);                     -- bresp
			f2h_BVALID                    : out   std_logic;                                        -- bvalid
			f2h_BREADY                    : in    std_logic                     := 'X';             -- bready
			f2h_ARID                      : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- arid
			f2h_ARADDR                    : in    std_logic_vector(31 downto 0) := (others => 'X'); -- araddr
			f2h_ARLEN                     : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- arlen
			f2h_ARSIZE                    : in    std_logic_vector(2 downto 0)  := (others => 'X'); -- arsize
			f2h_ARBURST                   : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- arburst
			f2h_ARLOCK                    : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- arlock
			f2h_ARCACHE                   : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- arcache
			f2h_ARPROT                    : in    std_logic_vector(2 downto 0)  := (others => 'X'); -- arprot
			f2h_ARVALID                   : in    std_logic                     := 'X';             -- arvalid
			f2h_ARREADY                   : out   std_logic;                                        -- arready
			f2h_ARUSER                    : in    std_logic_vector(4 downto 0)  := (others => 'X'); -- aruser
			f2h_RID                       : out   std_logic_vector(7 downto 0);                     -- rid
			f2h_RDATA                     : out   std_logic_vector(63 downto 0);                    -- rdata
			f2h_RRESP                     : out   std_logic_vector(1 downto 0);                     -- rresp
			f2h_RLAST                     : out   std_logic;                                        -- rlast
			f2h_RVALID                    : out   std_logic;                                        -- rvalid
			f2h_RREADY                    : in    std_logic                     := 'X';             -- rready
			h2f_lw_axi_clk                : in    std_logic                     := 'X';             -- clk
			h2f_lw_AWID                   : out   std_logic_vector(11 downto 0);                    -- awid
			h2f_lw_AWADDR                 : out   std_logic_vector(20 downto 0);                    -- awaddr
			h2f_lw_AWLEN                  : out   std_logic_vector(3 downto 0);                     -- awlen
			h2f_lw_AWSIZE                 : out   std_logic_vector(2 downto 0);                     -- awsize
			h2f_lw_AWBURST                : out   std_logic_vector(1 downto 0);                     -- awburst
			h2f_lw_AWLOCK                 : out   std_logic_vector(1 downto 0);                     -- awlock
			h2f_lw_AWCACHE                : out   std_logic_vector(3 downto 0);                     -- awcache
			h2f_lw_AWPROT                 : out   std_logic_vector(2 downto 0);                     -- awprot
			h2f_lw_AWVALID                : out   std_logic;                                        -- awvalid
			h2f_lw_AWREADY                : in    std_logic                     := 'X';             -- awready
			h2f_lw_WID                    : out   std_logic_vector(11 downto 0);                    -- wid
			h2f_lw_WDATA                  : out   std_logic_vector(31 downto 0);                    -- wdata
			h2f_lw_WSTRB                  : out   std_logic_vector(3 downto 0);                     -- wstrb
			h2f_lw_WLAST                  : out   std_logic;                                        -- wlast
			h2f_lw_WVALID                 : out   std_logic;                                        -- wvalid
			h2f_lw_WREADY                 : in    std_logic                     := 'X';             -- wready
			h2f_lw_BID                    : in    std_logic_vector(11 downto 0) := (others => 'X'); -- bid
			h2f_lw_BRESP                  : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- bresp
			h2f_lw_BVALID                 : in    std_logic                     := 'X';             -- bvalid
			h2f_lw_BREADY                 : out   std_logic;                                        -- bready
			h2f_lw_ARID                   : out   std_logic_vector(11 downto 0);                    -- arid
			h2f_lw_ARADDR                 : out   std_logic_vector(20 downto 0);                    -- araddr
			h2f_lw_ARLEN                  : out   std_logic_vector(3 downto 0);                     -- arlen
			h2f_lw_ARSIZE                 : out   std_logic_vector(2 downto 0);                     -- arsize
			h2f_lw_ARBURST                : out   std_logic_vector(1 downto 0);                     -- arburst
			h2f_lw_ARLOCK                 : out   std_logic_vector(1 downto 0);                     -- arlock
			h2f_lw_ARCACHE                : out   std_logic_vector(3 downto 0);                     -- arcache
			h2f_lw_ARPROT                 : out   std_logic_vector(2 downto 0);                     -- arprot
			h2f_lw_ARVALID                : out   std_logic;                                        -- arvalid
			h2f_lw_ARREADY                : in    std_logic                     := 'X';             -- arready
			h2f_lw_RID                    : in    std_logic_vector(11 downto 0) := (others => 'X'); -- rid
			h2f_lw_RDATA                  : in    std_logic_vector(31 downto 0) := (others => 'X'); -- rdata
			h2f_lw_RRESP                  : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- rresp
			h2f_lw_RLAST                  : in    std_logic                     := 'X';             -- rlast
			h2f_lw_RVALID                 : in    std_logic                     := 'X';             -- rvalid
			h2f_lw_RREADY                 : out   std_logic;                                        -- rready
			f2h_irq_p0                    : in    std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			f2h_irq_p1                    : in    std_logic_vector(31 downto 0) := (others => 'X')  -- irq
		);
	end component Computer_System_ARM_A9_HPS;

	component Computer_System_FPGA_Boot_SRAM is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(7 downto 0);                     -- readdata
			writedata  : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X'              -- reset_req
		);
	end component Computer_System_FPGA_Boot_SRAM;

	component Computer_System_JTAG_UART_for_ARM_0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component Computer_System_JTAG_UART_for_ARM_0;

	component Computer_System_JTAG_to_FPGA_Bridge is
		generic (
			USE_PLI     : integer := 0;
			PLI_PORT    : integer := 50000;
			FIFO_DEPTHS : integer := 2
		);
		port (
			clk_clk              : in  std_logic                     := 'X';             -- clk
			clk_reset_reset      : in  std_logic                     := 'X';             -- reset
			master_address       : out std_logic_vector(31 downto 0);                    -- address
			master_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			master_read          : out std_logic;                                        -- read
			master_write         : out std_logic;                                        -- write
			master_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			master_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			master_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			master_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			master_reset_reset   : out std_logic                                         -- reset
		);
	end component Computer_System_JTAG_to_FPGA_Bridge;

	component Computer_System_SysID is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component Computer_System_SysID;

	component Computer_System_System_PLL is
		port (
			ref_clk_clk        : in  std_logic := 'X'; -- clk
			ref_reset_reset    : in  std_logic := 'X'; -- reset
			sys_clk_clk        : out std_logic;        -- clk
			sdram_clk_clk      : out std_logic;        -- clk
			reset_source_reset : out std_logic         -- reset
		);
	end component Computer_System_System_PLL;

	component Computer_System_mm_interconnect_0 is
		port (
			ARM_A9_HPS_h2f_axi_master_awid                                        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- awid
			ARM_A9_HPS_h2f_axi_master_awaddr                                      : in  std_logic_vector(29 downto 0) := (others => 'X'); -- awaddr
			ARM_A9_HPS_h2f_axi_master_awlen                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awlen
			ARM_A9_HPS_h2f_axi_master_awsize                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awsize
			ARM_A9_HPS_h2f_axi_master_awburst                                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awburst
			ARM_A9_HPS_h2f_axi_master_awlock                                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awlock
			ARM_A9_HPS_h2f_axi_master_awcache                                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awcache
			ARM_A9_HPS_h2f_axi_master_awprot                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awprot
			ARM_A9_HPS_h2f_axi_master_awvalid                                     : in  std_logic                     := 'X';             -- awvalid
			ARM_A9_HPS_h2f_axi_master_awready                                     : out std_logic;                                        -- awready
			ARM_A9_HPS_h2f_axi_master_wid                                         : in  std_logic_vector(11 downto 0) := (others => 'X'); -- wid
			ARM_A9_HPS_h2f_axi_master_wdata                                       : in  std_logic_vector(63 downto 0) := (others => 'X'); -- wdata
			ARM_A9_HPS_h2f_axi_master_wstrb                                       : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- wstrb
			ARM_A9_HPS_h2f_axi_master_wlast                                       : in  std_logic                     := 'X';             -- wlast
			ARM_A9_HPS_h2f_axi_master_wvalid                                      : in  std_logic                     := 'X';             -- wvalid
			ARM_A9_HPS_h2f_axi_master_wready                                      : out std_logic;                                        -- wready
			ARM_A9_HPS_h2f_axi_master_bid                                         : out std_logic_vector(11 downto 0);                    -- bid
			ARM_A9_HPS_h2f_axi_master_bresp                                       : out std_logic_vector(1 downto 0);                     -- bresp
			ARM_A9_HPS_h2f_axi_master_bvalid                                      : out std_logic;                                        -- bvalid
			ARM_A9_HPS_h2f_axi_master_bready                                      : in  std_logic                     := 'X';             -- bready
			ARM_A9_HPS_h2f_axi_master_arid                                        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- arid
			ARM_A9_HPS_h2f_axi_master_araddr                                      : in  std_logic_vector(29 downto 0) := (others => 'X'); -- araddr
			ARM_A9_HPS_h2f_axi_master_arlen                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arlen
			ARM_A9_HPS_h2f_axi_master_arsize                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arsize
			ARM_A9_HPS_h2f_axi_master_arburst                                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arburst
			ARM_A9_HPS_h2f_axi_master_arlock                                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arlock
			ARM_A9_HPS_h2f_axi_master_arcache                                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arcache
			ARM_A9_HPS_h2f_axi_master_arprot                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arprot
			ARM_A9_HPS_h2f_axi_master_arvalid                                     : in  std_logic                     := 'X';             -- arvalid
			ARM_A9_HPS_h2f_axi_master_arready                                     : out std_logic;                                        -- arready
			ARM_A9_HPS_h2f_axi_master_rid                                         : out std_logic_vector(11 downto 0);                    -- rid
			ARM_A9_HPS_h2f_axi_master_rdata                                       : out std_logic_vector(63 downto 0);                    -- rdata
			ARM_A9_HPS_h2f_axi_master_rresp                                       : out std_logic_vector(1 downto 0);                     -- rresp
			ARM_A9_HPS_h2f_axi_master_rlast                                       : out std_logic;                                        -- rlast
			ARM_A9_HPS_h2f_axi_master_rvalid                                      : out std_logic;                                        -- rvalid
			ARM_A9_HPS_h2f_axi_master_rready                                      : in  std_logic                     := 'X';             -- rready
			ARM_A9_HPS_h2f_lw_axi_master_awid                                     : in  std_logic_vector(11 downto 0) := (others => 'X'); -- awid
			ARM_A9_HPS_h2f_lw_axi_master_awaddr                                   : in  std_logic_vector(20 downto 0) := (others => 'X'); -- awaddr
			ARM_A9_HPS_h2f_lw_axi_master_awlen                                    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awlen
			ARM_A9_HPS_h2f_lw_axi_master_awsize                                   : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awsize
			ARM_A9_HPS_h2f_lw_axi_master_awburst                                  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awburst
			ARM_A9_HPS_h2f_lw_axi_master_awlock                                   : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awlock
			ARM_A9_HPS_h2f_lw_axi_master_awcache                                  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awcache
			ARM_A9_HPS_h2f_lw_axi_master_awprot                                   : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awprot
			ARM_A9_HPS_h2f_lw_axi_master_awvalid                                  : in  std_logic                     := 'X';             -- awvalid
			ARM_A9_HPS_h2f_lw_axi_master_awready                                  : out std_logic;                                        -- awready
			ARM_A9_HPS_h2f_lw_axi_master_wid                                      : in  std_logic_vector(11 downto 0) := (others => 'X'); -- wid
			ARM_A9_HPS_h2f_lw_axi_master_wdata                                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wdata
			ARM_A9_HPS_h2f_lw_axi_master_wstrb                                    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- wstrb
			ARM_A9_HPS_h2f_lw_axi_master_wlast                                    : in  std_logic                     := 'X';             -- wlast
			ARM_A9_HPS_h2f_lw_axi_master_wvalid                                   : in  std_logic                     := 'X';             -- wvalid
			ARM_A9_HPS_h2f_lw_axi_master_wready                                   : out std_logic;                                        -- wready
			ARM_A9_HPS_h2f_lw_axi_master_bid                                      : out std_logic_vector(11 downto 0);                    -- bid
			ARM_A9_HPS_h2f_lw_axi_master_bresp                                    : out std_logic_vector(1 downto 0);                     -- bresp
			ARM_A9_HPS_h2f_lw_axi_master_bvalid                                   : out std_logic;                                        -- bvalid
			ARM_A9_HPS_h2f_lw_axi_master_bready                                   : in  std_logic                     := 'X';             -- bready
			ARM_A9_HPS_h2f_lw_axi_master_arid                                     : in  std_logic_vector(11 downto 0) := (others => 'X'); -- arid
			ARM_A9_HPS_h2f_lw_axi_master_araddr                                   : in  std_logic_vector(20 downto 0) := (others => 'X'); -- araddr
			ARM_A9_HPS_h2f_lw_axi_master_arlen                                    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arlen
			ARM_A9_HPS_h2f_lw_axi_master_arsize                                   : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arsize
			ARM_A9_HPS_h2f_lw_axi_master_arburst                                  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arburst
			ARM_A9_HPS_h2f_lw_axi_master_arlock                                   : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arlock
			ARM_A9_HPS_h2f_lw_axi_master_arcache                                  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arcache
			ARM_A9_HPS_h2f_lw_axi_master_arprot                                   : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arprot
			ARM_A9_HPS_h2f_lw_axi_master_arvalid                                  : in  std_logic                     := 'X';             -- arvalid
			ARM_A9_HPS_h2f_lw_axi_master_arready                                  : out std_logic;                                        -- arready
			ARM_A9_HPS_h2f_lw_axi_master_rid                                      : out std_logic_vector(11 downto 0);                    -- rid
			ARM_A9_HPS_h2f_lw_axi_master_rdata                                    : out std_logic_vector(31 downto 0);                    -- rdata
			ARM_A9_HPS_h2f_lw_axi_master_rresp                                    : out std_logic_vector(1 downto 0);                     -- rresp
			ARM_A9_HPS_h2f_lw_axi_master_rlast                                    : out std_logic;                                        -- rlast
			ARM_A9_HPS_h2f_lw_axi_master_rvalid                                   : out std_logic;                                        -- rvalid
			ARM_A9_HPS_h2f_lw_axi_master_rready                                   : in  std_logic                     := 'X';             -- rready
			System_PLL_sys_clk_clk                                                : in  std_logic                     := 'X';             -- clk
			ARM_A9_HPS_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			FPGA_Boot_SRAM_reset1_reset_bridge_in_reset_reset                     : in  std_logic                     := 'X';             -- reset
			JTAG_to_FPGA_Bridge_clk_reset_reset_bridge_in_reset_reset             : in  std_logic                     := 'X';             -- reset
			JTAG_to_FPGA_Bridge_master_address                                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			JTAG_to_FPGA_Bridge_master_waitrequest                                : out std_logic;                                        -- waitrequest
			JTAG_to_FPGA_Bridge_master_byteenable                                 : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			JTAG_to_FPGA_Bridge_master_read                                       : in  std_logic                     := 'X';             -- read
			JTAG_to_FPGA_Bridge_master_readdata                                   : out std_logic_vector(31 downto 0);                    -- readdata
			JTAG_to_FPGA_Bridge_master_readdatavalid                              : out std_logic;                                        -- readdatavalid
			JTAG_to_FPGA_Bridge_master_write                                      : in  std_logic                     := 'X';             -- write
			JTAG_to_FPGA_Bridge_master_writedata                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			FPGA_Boot_SRAM_s1_address                                             : out std_logic_vector(15 downto 0);                    -- address
			FPGA_Boot_SRAM_s1_write                                               : out std_logic;                                        -- write
			FPGA_Boot_SRAM_s1_readdata                                            : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			FPGA_Boot_SRAM_s1_writedata                                           : out std_logic_vector(7 downto 0);                     -- writedata
			FPGA_Boot_SRAM_s1_chipselect                                          : out std_logic;                                        -- chipselect
			FPGA_Boot_SRAM_s1_clken                                               : out std_logic;                                        -- clken
			JTAG_UART_for_ARM_0_avalon_jtag_slave_address                         : out std_logic_vector(0 downto 0);                     -- address
			JTAG_UART_for_ARM_0_avalon_jtag_slave_write                           : out std_logic;                                        -- write
			JTAG_UART_for_ARM_0_avalon_jtag_slave_read                            : out std_logic;                                        -- read
			JTAG_UART_for_ARM_0_avalon_jtag_slave_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			JTAG_UART_for_ARM_0_avalon_jtag_slave_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			JTAG_UART_for_ARM_0_avalon_jtag_slave_waitrequest                     : in  std_logic                     := 'X';             -- waitrequest
			JTAG_UART_for_ARM_0_avalon_jtag_slave_chipselect                      : out std_logic;                                        -- chipselect
			JTAG_UART_for_ARM_1_avalon_jtag_slave_address                         : out std_logic_vector(0 downto 0);                     -- address
			JTAG_UART_for_ARM_1_avalon_jtag_slave_write                           : out std_logic;                                        -- write
			JTAG_UART_for_ARM_1_avalon_jtag_slave_read                            : out std_logic;                                        -- read
			JTAG_UART_for_ARM_1_avalon_jtag_slave_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			JTAG_UART_for_ARM_1_avalon_jtag_slave_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			JTAG_UART_for_ARM_1_avalon_jtag_slave_waitrequest                     : in  std_logic                     := 'X';             -- waitrequest
			JTAG_UART_for_ARM_1_avalon_jtag_slave_chipselect                      : out std_logic;                                        -- chipselect
			SysID_control_slave_address                                           : out std_logic_vector(0 downto 0);                     -- address
			SysID_control_slave_readdata                                          : in  std_logic_vector(31 downto 0) := (others => 'X')  -- readdata
		);
	end component Computer_System_mm_interconnect_0;

	component Computer_System_mm_interconnect_1 is
		port (
			ARM_A9_HPS_f2h_axi_slave_awid                                          : out std_logic_vector(7 downto 0);                     -- awid
			ARM_A9_HPS_f2h_axi_slave_awaddr                                        : out std_logic_vector(31 downto 0);                    -- awaddr
			ARM_A9_HPS_f2h_axi_slave_awlen                                         : out std_logic_vector(3 downto 0);                     -- awlen
			ARM_A9_HPS_f2h_axi_slave_awsize                                        : out std_logic_vector(2 downto 0);                     -- awsize
			ARM_A9_HPS_f2h_axi_slave_awburst                                       : out std_logic_vector(1 downto 0);                     -- awburst
			ARM_A9_HPS_f2h_axi_slave_awlock                                        : out std_logic_vector(1 downto 0);                     -- awlock
			ARM_A9_HPS_f2h_axi_slave_awcache                                       : out std_logic_vector(3 downto 0);                     -- awcache
			ARM_A9_HPS_f2h_axi_slave_awprot                                        : out std_logic_vector(2 downto 0);                     -- awprot
			ARM_A9_HPS_f2h_axi_slave_awuser                                        : out std_logic_vector(4 downto 0);                     -- awuser
			ARM_A9_HPS_f2h_axi_slave_awvalid                                       : out std_logic;                                        -- awvalid
			ARM_A9_HPS_f2h_axi_slave_awready                                       : in  std_logic                     := 'X';             -- awready
			ARM_A9_HPS_f2h_axi_slave_wid                                           : out std_logic_vector(7 downto 0);                     -- wid
			ARM_A9_HPS_f2h_axi_slave_wdata                                         : out std_logic_vector(63 downto 0);                    -- wdata
			ARM_A9_HPS_f2h_axi_slave_wstrb                                         : out std_logic_vector(7 downto 0);                     -- wstrb
			ARM_A9_HPS_f2h_axi_slave_wlast                                         : out std_logic;                                        -- wlast
			ARM_A9_HPS_f2h_axi_slave_wvalid                                        : out std_logic;                                        -- wvalid
			ARM_A9_HPS_f2h_axi_slave_wready                                        : in  std_logic                     := 'X';             -- wready
			ARM_A9_HPS_f2h_axi_slave_bid                                           : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- bid
			ARM_A9_HPS_f2h_axi_slave_bresp                                         : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- bresp
			ARM_A9_HPS_f2h_axi_slave_bvalid                                        : in  std_logic                     := 'X';             -- bvalid
			ARM_A9_HPS_f2h_axi_slave_bready                                        : out std_logic;                                        -- bready
			ARM_A9_HPS_f2h_axi_slave_arid                                          : out std_logic_vector(7 downto 0);                     -- arid
			ARM_A9_HPS_f2h_axi_slave_araddr                                        : out std_logic_vector(31 downto 0);                    -- araddr
			ARM_A9_HPS_f2h_axi_slave_arlen                                         : out std_logic_vector(3 downto 0);                     -- arlen
			ARM_A9_HPS_f2h_axi_slave_arsize                                        : out std_logic_vector(2 downto 0);                     -- arsize
			ARM_A9_HPS_f2h_axi_slave_arburst                                       : out std_logic_vector(1 downto 0);                     -- arburst
			ARM_A9_HPS_f2h_axi_slave_arlock                                        : out std_logic_vector(1 downto 0);                     -- arlock
			ARM_A9_HPS_f2h_axi_slave_arcache                                       : out std_logic_vector(3 downto 0);                     -- arcache
			ARM_A9_HPS_f2h_axi_slave_arprot                                        : out std_logic_vector(2 downto 0);                     -- arprot
			ARM_A9_HPS_f2h_axi_slave_aruser                                        : out std_logic_vector(4 downto 0);                     -- aruser
			ARM_A9_HPS_f2h_axi_slave_arvalid                                       : out std_logic;                                        -- arvalid
			ARM_A9_HPS_f2h_axi_slave_arready                                       : in  std_logic                     := 'X';             -- arready
			ARM_A9_HPS_f2h_axi_slave_rid                                           : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- rid
			ARM_A9_HPS_f2h_axi_slave_rdata                                         : in  std_logic_vector(63 downto 0) := (others => 'X'); -- rdata
			ARM_A9_HPS_f2h_axi_slave_rresp                                         : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- rresp
			ARM_A9_HPS_f2h_axi_slave_rlast                                         : in  std_logic                     := 'X';             -- rlast
			ARM_A9_HPS_f2h_axi_slave_rvalid                                        : in  std_logic                     := 'X';             -- rvalid
			ARM_A9_HPS_f2h_axi_slave_rready                                        : out std_logic;                                        -- rready
			System_PLL_sys_clk_clk                                                 : in  std_logic                     := 'X';             -- clk
			ARM_A9_HPS_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset_reset  : in  std_logic                     := 'X';             -- reset
			JTAG_to_HPS_Bridge_clk_reset_reset_bridge_in_reset_reset               : in  std_logic                     := 'X';             -- reset
			JTAG_to_HPS_Bridge_master_translator_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			JTAG_to_HPS_Bridge_master_address                                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			JTAG_to_HPS_Bridge_master_waitrequest                                  : out std_logic;                                        -- waitrequest
			JTAG_to_HPS_Bridge_master_byteenable                                   : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			JTAG_to_HPS_Bridge_master_read                                         : in  std_logic                     := 'X';             -- read
			JTAG_to_HPS_Bridge_master_readdata                                     : out std_logic_vector(31 downto 0);                    -- readdata
			JTAG_to_HPS_Bridge_master_readdatavalid                                : out std_logic;                                        -- readdatavalid
			JTAG_to_HPS_Bridge_master_write                                        : in  std_logic                     := 'X';             -- write
			JTAG_to_HPS_Bridge_master_writedata                                    : in  std_logic_vector(31 downto 0) := (others => 'X')  -- writedata
		);
	end component Computer_System_mm_interconnect_1;

	component Computer_System_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component Computer_System_irq_mapper;

	component computer_system_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component computer_system_rst_controller;

	component computer_system_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component computer_system_rst_controller_001;

	signal arm_a9_hps_h2f_reset_reset                                              : std_logic;                     -- ARM_A9_HPS:h2f_rst_n -> [fpga_reset_reset_n, fpga_reset_reset_n:in]
	signal system_pll_sys_clk_clk                                                  : std_logic;                     -- System_PLL:sys_clk_clk -> [ARM_A9_HPS:f2h_axi_clk, ARM_A9_HPS:h2f_axi_clk, ARM_A9_HPS:h2f_lw_axi_clk, FPGA_Boot_SRAM:clk, JTAG_UART_for_ARM_0:clk, JTAG_UART_for_ARM_1:clk, JTAG_to_FPGA_Bridge:clk_clk, JTAG_to_HPS_Bridge:clk_clk, SysID:clock, mm_interconnect_0:System_PLL_sys_clk_clk, mm_interconnect_1:System_PLL_sys_clk_clk, rst_controller:clk, rst_controller_001:clk]
	signal system_pll_reset_source_reset                                           : std_logic;                     -- System_PLL:reset_source_reset -> [JTAG_to_FPGA_Bridge:clk_reset_reset, JTAG_to_HPS_Bridge:clk_reset_reset, rst_controller:reset_in0]
	signal arm_a9_hps_h2f_axi_master_awburst                                       : std_logic_vector(1 downto 0);  -- ARM_A9_HPS:h2f_AWBURST -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awburst
	signal arm_a9_hps_h2f_axi_master_arlen                                         : std_logic_vector(3 downto 0);  -- ARM_A9_HPS:h2f_ARLEN -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arlen
	signal arm_a9_hps_h2f_axi_master_wstrb                                         : std_logic_vector(7 downto 0);  -- ARM_A9_HPS:h2f_WSTRB -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_wstrb
	signal arm_a9_hps_h2f_axi_master_wready                                        : std_logic;                     -- mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_wready -> ARM_A9_HPS:h2f_WREADY
	signal arm_a9_hps_h2f_axi_master_rid                                           : std_logic_vector(11 downto 0); -- mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_rid -> ARM_A9_HPS:h2f_RID
	signal arm_a9_hps_h2f_axi_master_rready                                        : std_logic;                     -- ARM_A9_HPS:h2f_RREADY -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_rready
	signal arm_a9_hps_h2f_axi_master_awlen                                         : std_logic_vector(3 downto 0);  -- ARM_A9_HPS:h2f_AWLEN -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awlen
	signal arm_a9_hps_h2f_axi_master_wid                                           : std_logic_vector(11 downto 0); -- ARM_A9_HPS:h2f_WID -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_wid
	signal arm_a9_hps_h2f_axi_master_arcache                                       : std_logic_vector(3 downto 0);  -- ARM_A9_HPS:h2f_ARCACHE -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arcache
	signal arm_a9_hps_h2f_axi_master_wvalid                                        : std_logic;                     -- ARM_A9_HPS:h2f_WVALID -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_wvalid
	signal arm_a9_hps_h2f_axi_master_araddr                                        : std_logic_vector(29 downto 0); -- ARM_A9_HPS:h2f_ARADDR -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_araddr
	signal arm_a9_hps_h2f_axi_master_arprot                                        : std_logic_vector(2 downto 0);  -- ARM_A9_HPS:h2f_ARPROT -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arprot
	signal arm_a9_hps_h2f_axi_master_awprot                                        : std_logic_vector(2 downto 0);  -- ARM_A9_HPS:h2f_AWPROT -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awprot
	signal arm_a9_hps_h2f_axi_master_wdata                                         : std_logic_vector(63 downto 0); -- ARM_A9_HPS:h2f_WDATA -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_wdata
	signal arm_a9_hps_h2f_axi_master_arvalid                                       : std_logic;                     -- ARM_A9_HPS:h2f_ARVALID -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arvalid
	signal arm_a9_hps_h2f_axi_master_awcache                                       : std_logic_vector(3 downto 0);  -- ARM_A9_HPS:h2f_AWCACHE -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awcache
	signal arm_a9_hps_h2f_axi_master_arid                                          : std_logic_vector(11 downto 0); -- ARM_A9_HPS:h2f_ARID -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arid
	signal arm_a9_hps_h2f_axi_master_arlock                                        : std_logic_vector(1 downto 0);  -- ARM_A9_HPS:h2f_ARLOCK -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arlock
	signal arm_a9_hps_h2f_axi_master_awlock                                        : std_logic_vector(1 downto 0);  -- ARM_A9_HPS:h2f_AWLOCK -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awlock
	signal arm_a9_hps_h2f_axi_master_awaddr                                        : std_logic_vector(29 downto 0); -- ARM_A9_HPS:h2f_AWADDR -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awaddr
	signal arm_a9_hps_h2f_axi_master_bresp                                         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_bresp -> ARM_A9_HPS:h2f_BRESP
	signal arm_a9_hps_h2f_axi_master_arready                                       : std_logic;                     -- mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arready -> ARM_A9_HPS:h2f_ARREADY
	signal arm_a9_hps_h2f_axi_master_rdata                                         : std_logic_vector(63 downto 0); -- mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_rdata -> ARM_A9_HPS:h2f_RDATA
	signal arm_a9_hps_h2f_axi_master_awready                                       : std_logic;                     -- mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awready -> ARM_A9_HPS:h2f_AWREADY
	signal arm_a9_hps_h2f_axi_master_arburst                                       : std_logic_vector(1 downto 0);  -- ARM_A9_HPS:h2f_ARBURST -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arburst
	signal arm_a9_hps_h2f_axi_master_arsize                                        : std_logic_vector(2 downto 0);  -- ARM_A9_HPS:h2f_ARSIZE -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arsize
	signal arm_a9_hps_h2f_axi_master_bready                                        : std_logic;                     -- ARM_A9_HPS:h2f_BREADY -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_bready
	signal arm_a9_hps_h2f_axi_master_rlast                                         : std_logic;                     -- mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_rlast -> ARM_A9_HPS:h2f_RLAST
	signal arm_a9_hps_h2f_axi_master_wlast                                         : std_logic;                     -- ARM_A9_HPS:h2f_WLAST -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_wlast
	signal arm_a9_hps_h2f_axi_master_rresp                                         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_rresp -> ARM_A9_HPS:h2f_RRESP
	signal arm_a9_hps_h2f_axi_master_awid                                          : std_logic_vector(11 downto 0); -- ARM_A9_HPS:h2f_AWID -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awid
	signal arm_a9_hps_h2f_axi_master_bid                                           : std_logic_vector(11 downto 0); -- mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_bid -> ARM_A9_HPS:h2f_BID
	signal arm_a9_hps_h2f_axi_master_bvalid                                        : std_logic;                     -- mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_bvalid -> ARM_A9_HPS:h2f_BVALID
	signal arm_a9_hps_h2f_axi_master_awsize                                        : std_logic_vector(2 downto 0);  -- ARM_A9_HPS:h2f_AWSIZE -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awsize
	signal arm_a9_hps_h2f_axi_master_awvalid                                       : std_logic;                     -- ARM_A9_HPS:h2f_AWVALID -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awvalid
	signal arm_a9_hps_h2f_axi_master_rvalid                                        : std_logic;                     -- mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_rvalid -> ARM_A9_HPS:h2f_RVALID
	signal jtag_to_fpga_bridge_master_readdata                                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:JTAG_to_FPGA_Bridge_master_readdata -> JTAG_to_FPGA_Bridge:master_readdata
	signal jtag_to_fpga_bridge_master_waitrequest                                  : std_logic;                     -- mm_interconnect_0:JTAG_to_FPGA_Bridge_master_waitrequest -> JTAG_to_FPGA_Bridge:master_waitrequest
	signal jtag_to_fpga_bridge_master_address                                      : std_logic_vector(31 downto 0); -- JTAG_to_FPGA_Bridge:master_address -> mm_interconnect_0:JTAG_to_FPGA_Bridge_master_address
	signal jtag_to_fpga_bridge_master_read                                         : std_logic;                     -- JTAG_to_FPGA_Bridge:master_read -> mm_interconnect_0:JTAG_to_FPGA_Bridge_master_read
	signal jtag_to_fpga_bridge_master_byteenable                                   : std_logic_vector(3 downto 0);  -- JTAG_to_FPGA_Bridge:master_byteenable -> mm_interconnect_0:JTAG_to_FPGA_Bridge_master_byteenable
	signal jtag_to_fpga_bridge_master_readdatavalid                                : std_logic;                     -- mm_interconnect_0:JTAG_to_FPGA_Bridge_master_readdatavalid -> JTAG_to_FPGA_Bridge:master_readdatavalid
	signal jtag_to_fpga_bridge_master_write                                        : std_logic;                     -- JTAG_to_FPGA_Bridge:master_write -> mm_interconnect_0:JTAG_to_FPGA_Bridge_master_write
	signal jtag_to_fpga_bridge_master_writedata                                    : std_logic_vector(31 downto 0); -- JTAG_to_FPGA_Bridge:master_writedata -> mm_interconnect_0:JTAG_to_FPGA_Bridge_master_writedata
	signal arm_a9_hps_h2f_lw_axi_master_awburst                                    : std_logic_vector(1 downto 0);  -- ARM_A9_HPS:h2f_lw_AWBURST -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awburst
	signal arm_a9_hps_h2f_lw_axi_master_arlen                                      : std_logic_vector(3 downto 0);  -- ARM_A9_HPS:h2f_lw_ARLEN -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arlen
	signal arm_a9_hps_h2f_lw_axi_master_wstrb                                      : std_logic_vector(3 downto 0);  -- ARM_A9_HPS:h2f_lw_WSTRB -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_wstrb
	signal arm_a9_hps_h2f_lw_axi_master_wready                                     : std_logic;                     -- mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_wready -> ARM_A9_HPS:h2f_lw_WREADY
	signal arm_a9_hps_h2f_lw_axi_master_rid                                        : std_logic_vector(11 downto 0); -- mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_rid -> ARM_A9_HPS:h2f_lw_RID
	signal arm_a9_hps_h2f_lw_axi_master_rready                                     : std_logic;                     -- ARM_A9_HPS:h2f_lw_RREADY -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_rready
	signal arm_a9_hps_h2f_lw_axi_master_awlen                                      : std_logic_vector(3 downto 0);  -- ARM_A9_HPS:h2f_lw_AWLEN -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awlen
	signal arm_a9_hps_h2f_lw_axi_master_wid                                        : std_logic_vector(11 downto 0); -- ARM_A9_HPS:h2f_lw_WID -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_wid
	signal arm_a9_hps_h2f_lw_axi_master_arcache                                    : std_logic_vector(3 downto 0);  -- ARM_A9_HPS:h2f_lw_ARCACHE -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arcache
	signal arm_a9_hps_h2f_lw_axi_master_wvalid                                     : std_logic;                     -- ARM_A9_HPS:h2f_lw_WVALID -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_wvalid
	signal arm_a9_hps_h2f_lw_axi_master_araddr                                     : std_logic_vector(20 downto 0); -- ARM_A9_HPS:h2f_lw_ARADDR -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_araddr
	signal arm_a9_hps_h2f_lw_axi_master_arprot                                     : std_logic_vector(2 downto 0);  -- ARM_A9_HPS:h2f_lw_ARPROT -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arprot
	signal arm_a9_hps_h2f_lw_axi_master_awprot                                     : std_logic_vector(2 downto 0);  -- ARM_A9_HPS:h2f_lw_AWPROT -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awprot
	signal arm_a9_hps_h2f_lw_axi_master_wdata                                      : std_logic_vector(31 downto 0); -- ARM_A9_HPS:h2f_lw_WDATA -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_wdata
	signal arm_a9_hps_h2f_lw_axi_master_arvalid                                    : std_logic;                     -- ARM_A9_HPS:h2f_lw_ARVALID -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arvalid
	signal arm_a9_hps_h2f_lw_axi_master_awcache                                    : std_logic_vector(3 downto 0);  -- ARM_A9_HPS:h2f_lw_AWCACHE -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awcache
	signal arm_a9_hps_h2f_lw_axi_master_arid                                       : std_logic_vector(11 downto 0); -- ARM_A9_HPS:h2f_lw_ARID -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arid
	signal arm_a9_hps_h2f_lw_axi_master_arlock                                     : std_logic_vector(1 downto 0);  -- ARM_A9_HPS:h2f_lw_ARLOCK -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arlock
	signal arm_a9_hps_h2f_lw_axi_master_awlock                                     : std_logic_vector(1 downto 0);  -- ARM_A9_HPS:h2f_lw_AWLOCK -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awlock
	signal arm_a9_hps_h2f_lw_axi_master_awaddr                                     : std_logic_vector(20 downto 0); -- ARM_A9_HPS:h2f_lw_AWADDR -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awaddr
	signal arm_a9_hps_h2f_lw_axi_master_bresp                                      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_bresp -> ARM_A9_HPS:h2f_lw_BRESP
	signal arm_a9_hps_h2f_lw_axi_master_arready                                    : std_logic;                     -- mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arready -> ARM_A9_HPS:h2f_lw_ARREADY
	signal arm_a9_hps_h2f_lw_axi_master_rdata                                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_rdata -> ARM_A9_HPS:h2f_lw_RDATA
	signal arm_a9_hps_h2f_lw_axi_master_awready                                    : std_logic;                     -- mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awready -> ARM_A9_HPS:h2f_lw_AWREADY
	signal arm_a9_hps_h2f_lw_axi_master_arburst                                    : std_logic_vector(1 downto 0);  -- ARM_A9_HPS:h2f_lw_ARBURST -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arburst
	signal arm_a9_hps_h2f_lw_axi_master_arsize                                     : std_logic_vector(2 downto 0);  -- ARM_A9_HPS:h2f_lw_ARSIZE -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_arsize
	signal arm_a9_hps_h2f_lw_axi_master_bready                                     : std_logic;                     -- ARM_A9_HPS:h2f_lw_BREADY -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_bready
	signal arm_a9_hps_h2f_lw_axi_master_rlast                                      : std_logic;                     -- mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_rlast -> ARM_A9_HPS:h2f_lw_RLAST
	signal arm_a9_hps_h2f_lw_axi_master_wlast                                      : std_logic;                     -- ARM_A9_HPS:h2f_lw_WLAST -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_wlast
	signal arm_a9_hps_h2f_lw_axi_master_rresp                                      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_rresp -> ARM_A9_HPS:h2f_lw_RRESP
	signal arm_a9_hps_h2f_lw_axi_master_awid                                       : std_logic_vector(11 downto 0); -- ARM_A9_HPS:h2f_lw_AWID -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awid
	signal arm_a9_hps_h2f_lw_axi_master_bid                                        : std_logic_vector(11 downto 0); -- mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_bid -> ARM_A9_HPS:h2f_lw_BID
	signal arm_a9_hps_h2f_lw_axi_master_bvalid                                     : std_logic;                     -- mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_bvalid -> ARM_A9_HPS:h2f_lw_BVALID
	signal arm_a9_hps_h2f_lw_axi_master_awsize                                     : std_logic_vector(2 downto 0);  -- ARM_A9_HPS:h2f_lw_AWSIZE -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awsize
	signal arm_a9_hps_h2f_lw_axi_master_awvalid                                    : std_logic;                     -- ARM_A9_HPS:h2f_lw_AWVALID -> mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_awvalid
	signal arm_a9_hps_h2f_lw_axi_master_rvalid                                     : std_logic;                     -- mm_interconnect_0:ARM_A9_HPS_h2f_lw_axi_master_rvalid -> ARM_A9_HPS:h2f_lw_RVALID
	signal mm_interconnect_0_fpga_boot_sram_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:FPGA_Boot_SRAM_s1_chipselect -> FPGA_Boot_SRAM:chipselect
	signal mm_interconnect_0_fpga_boot_sram_s1_readdata                            : std_logic_vector(7 downto 0);  -- FPGA_Boot_SRAM:readdata -> mm_interconnect_0:FPGA_Boot_SRAM_s1_readdata
	signal mm_interconnect_0_fpga_boot_sram_s1_address                             : std_logic_vector(15 downto 0); -- mm_interconnect_0:FPGA_Boot_SRAM_s1_address -> FPGA_Boot_SRAM:address
	signal mm_interconnect_0_fpga_boot_sram_s1_write                               : std_logic;                     -- mm_interconnect_0:FPGA_Boot_SRAM_s1_write -> FPGA_Boot_SRAM:write
	signal mm_interconnect_0_fpga_boot_sram_s1_writedata                           : std_logic_vector(7 downto 0);  -- mm_interconnect_0:FPGA_Boot_SRAM_s1_writedata -> FPGA_Boot_SRAM:writedata
	signal mm_interconnect_0_fpga_boot_sram_s1_clken                               : std_logic;                     -- mm_interconnect_0:FPGA_Boot_SRAM_s1_clken -> FPGA_Boot_SRAM:clken
	signal mm_interconnect_0_sysid_control_slave_readdata                          : std_logic_vector(31 downto 0); -- SysID:readdata -> mm_interconnect_0:SysID_control_slave_readdata
	signal mm_interconnect_0_sysid_control_slave_address                           : std_logic_vector(0 downto 0);  -- mm_interconnect_0:SysID_control_slave_address -> SysID:address
	signal mm_interconnect_0_jtag_uart_for_arm_0_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:JTAG_UART_for_ARM_0_avalon_jtag_slave_chipselect -> JTAG_UART_for_ARM_0:av_chipselect
	signal mm_interconnect_0_jtag_uart_for_arm_0_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- JTAG_UART_for_ARM_0:av_readdata -> mm_interconnect_0:JTAG_UART_for_ARM_0_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_for_arm_0_avalon_jtag_slave_waitrequest     : std_logic;                     -- JTAG_UART_for_ARM_0:av_waitrequest -> mm_interconnect_0:JTAG_UART_for_ARM_0_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_for_arm_0_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:JTAG_UART_for_ARM_0_avalon_jtag_slave_address -> JTAG_UART_for_ARM_0:av_address
	signal mm_interconnect_0_jtag_uart_for_arm_0_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:JTAG_UART_for_ARM_0_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_for_arm_0_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_for_arm_0_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:JTAG_UART_for_ARM_0_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_for_arm_0_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_for_arm_0_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:JTAG_UART_for_ARM_0_avalon_jtag_slave_writedata -> JTAG_UART_for_ARM_0:av_writedata
	signal mm_interconnect_0_jtag_uart_for_arm_1_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:JTAG_UART_for_ARM_1_avalon_jtag_slave_chipselect -> JTAG_UART_for_ARM_1:av_chipselect
	signal mm_interconnect_0_jtag_uart_for_arm_1_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- JTAG_UART_for_ARM_1:av_readdata -> mm_interconnect_0:JTAG_UART_for_ARM_1_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_for_arm_1_avalon_jtag_slave_waitrequest     : std_logic;                     -- JTAG_UART_for_ARM_1:av_waitrequest -> mm_interconnect_0:JTAG_UART_for_ARM_1_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_for_arm_1_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:JTAG_UART_for_ARM_1_avalon_jtag_slave_address -> JTAG_UART_for_ARM_1:av_address
	signal mm_interconnect_0_jtag_uart_for_arm_1_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:JTAG_UART_for_ARM_1_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_for_arm_1_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_for_arm_1_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:JTAG_UART_for_ARM_1_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_for_arm_1_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_for_arm_1_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:JTAG_UART_for_ARM_1_avalon_jtag_slave_writedata -> JTAG_UART_for_ARM_1:av_writedata
	signal jtag_to_hps_bridge_master_readdata                                      : std_logic_vector(31 downto 0); -- mm_interconnect_1:JTAG_to_HPS_Bridge_master_readdata -> JTAG_to_HPS_Bridge:master_readdata
	signal jtag_to_hps_bridge_master_waitrequest                                   : std_logic;                     -- mm_interconnect_1:JTAG_to_HPS_Bridge_master_waitrequest -> JTAG_to_HPS_Bridge:master_waitrequest
	signal jtag_to_hps_bridge_master_address                                       : std_logic_vector(31 downto 0); -- JTAG_to_HPS_Bridge:master_address -> mm_interconnect_1:JTAG_to_HPS_Bridge_master_address
	signal jtag_to_hps_bridge_master_read                                          : std_logic;                     -- JTAG_to_HPS_Bridge:master_read -> mm_interconnect_1:JTAG_to_HPS_Bridge_master_read
	signal jtag_to_hps_bridge_master_byteenable                                    : std_logic_vector(3 downto 0);  -- JTAG_to_HPS_Bridge:master_byteenable -> mm_interconnect_1:JTAG_to_HPS_Bridge_master_byteenable
	signal jtag_to_hps_bridge_master_readdatavalid                                 : std_logic;                     -- mm_interconnect_1:JTAG_to_HPS_Bridge_master_readdatavalid -> JTAG_to_HPS_Bridge:master_readdatavalid
	signal jtag_to_hps_bridge_master_write                                         : std_logic;                     -- JTAG_to_HPS_Bridge:master_write -> mm_interconnect_1:JTAG_to_HPS_Bridge_master_write
	signal jtag_to_hps_bridge_master_writedata                                     : std_logic_vector(31 downto 0); -- JTAG_to_HPS_Bridge:master_writedata -> mm_interconnect_1:JTAG_to_HPS_Bridge_master_writedata
	signal mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awburst                      : std_logic_vector(1 downto 0);  -- mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_awburst -> ARM_A9_HPS:f2h_AWBURST
	signal mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awuser                       : std_logic_vector(4 downto 0);  -- mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_awuser -> ARM_A9_HPS:f2h_AWUSER
	signal mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arlen                        : std_logic_vector(3 downto 0);  -- mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_arlen -> ARM_A9_HPS:f2h_ARLEN
	signal mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wstrb                        : std_logic_vector(7 downto 0);  -- mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_wstrb -> ARM_A9_HPS:f2h_WSTRB
	signal mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wready                       : std_logic;                     -- ARM_A9_HPS:f2h_WREADY -> mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_wready
	signal mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rid                          : std_logic_vector(7 downto 0);  -- ARM_A9_HPS:f2h_RID -> mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_rid
	signal mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rready                       : std_logic;                     -- mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_rready -> ARM_A9_HPS:f2h_RREADY
	signal mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awlen                        : std_logic_vector(3 downto 0);  -- mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_awlen -> ARM_A9_HPS:f2h_AWLEN
	signal mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wid                          : std_logic_vector(7 downto 0);  -- mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_wid -> ARM_A9_HPS:f2h_WID
	signal mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arcache                      : std_logic_vector(3 downto 0);  -- mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_arcache -> ARM_A9_HPS:f2h_ARCACHE
	signal mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wvalid                       : std_logic;                     -- mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_wvalid -> ARM_A9_HPS:f2h_WVALID
	signal mm_interconnect_1_arm_a9_hps_f2h_axi_slave_araddr                       : std_logic_vector(31 downto 0); -- mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_araddr -> ARM_A9_HPS:f2h_ARADDR
	signal mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arprot                       : std_logic_vector(2 downto 0);  -- mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_arprot -> ARM_A9_HPS:f2h_ARPROT
	signal mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awprot                       : std_logic_vector(2 downto 0);  -- mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_awprot -> ARM_A9_HPS:f2h_AWPROT
	signal mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wdata                        : std_logic_vector(63 downto 0); -- mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_wdata -> ARM_A9_HPS:f2h_WDATA
	signal mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arvalid                      : std_logic;                     -- mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_arvalid -> ARM_A9_HPS:f2h_ARVALID
	signal mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awcache                      : std_logic_vector(3 downto 0);  -- mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_awcache -> ARM_A9_HPS:f2h_AWCACHE
	signal mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arid                         : std_logic_vector(7 downto 0);  -- mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_arid -> ARM_A9_HPS:f2h_ARID
	signal mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arlock                       : std_logic_vector(1 downto 0);  -- mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_arlock -> ARM_A9_HPS:f2h_ARLOCK
	signal mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awlock                       : std_logic_vector(1 downto 0);  -- mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_awlock -> ARM_A9_HPS:f2h_AWLOCK
	signal mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awaddr                       : std_logic_vector(31 downto 0); -- mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_awaddr -> ARM_A9_HPS:f2h_AWADDR
	signal mm_interconnect_1_arm_a9_hps_f2h_axi_slave_bresp                        : std_logic_vector(1 downto 0);  -- ARM_A9_HPS:f2h_BRESP -> mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_bresp
	signal mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arready                      : std_logic;                     -- ARM_A9_HPS:f2h_ARREADY -> mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_arready
	signal mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rdata                        : std_logic_vector(63 downto 0); -- ARM_A9_HPS:f2h_RDATA -> mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_rdata
	signal mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awready                      : std_logic;                     -- ARM_A9_HPS:f2h_AWREADY -> mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_awready
	signal mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arburst                      : std_logic_vector(1 downto 0);  -- mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_arburst -> ARM_A9_HPS:f2h_ARBURST
	signal mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arsize                       : std_logic_vector(2 downto 0);  -- mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_arsize -> ARM_A9_HPS:f2h_ARSIZE
	signal mm_interconnect_1_arm_a9_hps_f2h_axi_slave_bready                       : std_logic;                     -- mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_bready -> ARM_A9_HPS:f2h_BREADY
	signal mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rlast                        : std_logic;                     -- ARM_A9_HPS:f2h_RLAST -> mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_rlast
	signal mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wlast                        : std_logic;                     -- mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_wlast -> ARM_A9_HPS:f2h_WLAST
	signal mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rresp                        : std_logic_vector(1 downto 0);  -- ARM_A9_HPS:f2h_RRESP -> mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_rresp
	signal mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awid                         : std_logic_vector(7 downto 0);  -- mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_awid -> ARM_A9_HPS:f2h_AWID
	signal mm_interconnect_1_arm_a9_hps_f2h_axi_slave_bid                          : std_logic_vector(7 downto 0);  -- ARM_A9_HPS:f2h_BID -> mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_bid
	signal mm_interconnect_1_arm_a9_hps_f2h_axi_slave_bvalid                       : std_logic;                     -- ARM_A9_HPS:f2h_BVALID -> mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_bvalid
	signal mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awsize                       : std_logic_vector(2 downto 0);  -- mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_awsize -> ARM_A9_HPS:f2h_AWSIZE
	signal mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awvalid                      : std_logic;                     -- mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_awvalid -> ARM_A9_HPS:f2h_AWVALID
	signal mm_interconnect_1_arm_a9_hps_f2h_axi_slave_aruser                       : std_logic_vector(4 downto 0);  -- mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_aruser -> ARM_A9_HPS:f2h_ARUSER
	signal mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rvalid                       : std_logic;                     -- ARM_A9_HPS:f2h_RVALID -> mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_rvalid
	signal irq_mapper_receiver0_irq                                                : std_logic;                     -- JTAG_UART_for_ARM_0:av_irq -> irq_mapper:receiver0_irq
	signal arm_a9_hps_f2h_irq0_irq                                                 : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> ARM_A9_HPS:f2h_irq_p0
	signal irq_mapper_001_receiver0_irq                                            : std_logic;                     -- JTAG_UART_for_ARM_1:av_irq -> irq_mapper_001:receiver0_irq
	signal arm_a9_hps_f2h_irq1_irq                                                 : std_logic_vector(31 downto 0); -- irq_mapper_001:sender_irq -> ARM_A9_HPS:f2h_irq_p1
	signal rst_controller_reset_out_reset                                          : std_logic;                     -- rst_controller:reset_out -> [FPGA_Boot_SRAM:reset, mm_interconnect_0:FPGA_Boot_SRAM_reset1_reset_bridge_in_reset_reset, mm_interconnect_0:JTAG_to_FPGA_Bridge_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_1:JTAG_to_HPS_Bridge_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_1:JTAG_to_HPS_Bridge_master_translator_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                                      : std_logic;                     -- rst_controller:reset_req -> [FPGA_Boot_SRAM:reset_req, rst_translator:reset_req_in]
	signal rst_controller_001_reset_out_reset                                      : std_logic;                     -- rst_controller_001:reset_out -> [mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_1:ARM_A9_HPS_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset_reset]
	signal fpga_reset_reset_n_ports_inv                                            : std_logic;                     -- fpga_reset_reset_n:inv -> rst_controller_001:reset_in0
	signal mm_interconnect_0_jtag_uart_for_arm_0_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_for_arm_0_avalon_jtag_slave_read:inv -> JTAG_UART_for_ARM_0:av_read_n
	signal mm_interconnect_0_jtag_uart_for_arm_0_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_uart_for_arm_0_avalon_jtag_slave_write:inv -> JTAG_UART_for_ARM_0:av_write_n
	signal mm_interconnect_0_jtag_uart_for_arm_1_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_for_arm_1_avalon_jtag_slave_read:inv -> JTAG_UART_for_ARM_1:av_read_n
	signal mm_interconnect_0_jtag_uart_for_arm_1_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_uart_for_arm_1_avalon_jtag_slave_write:inv -> JTAG_UART_for_ARM_1:av_write_n
	signal rst_controller_reset_out_reset_ports_inv                                : std_logic;                     -- rst_controller_reset_out_reset:inv -> [JTAG_UART_for_ARM_0:rst_n, JTAG_UART_for_ARM_1:rst_n, SysID:reset_n]

begin

	arm_a9_hps : component Computer_System_ARM_A9_HPS
		generic map (
			F2S_Width => 2,
			S2F_Width => 2
		)
		port map (
			h2f_loan_in                   => h2f_loan_io_in,                                     --        h2f_loan_io.in
			h2f_loan_out                  => h2f_loan_io_out,                                    --                   .out
			h2f_loan_oe                   => h2f_loan_io_oe,                                     --                   .oe
			f2h_boot_from_fpga_ready      => f2h_bootflags_boot_from_fpga_ready,                 -- f2h_boot_from_fpga.boot_from_fpga_ready
			f2h_boot_from_fpga_on_failure => f2h_bootflags_boot_from_fpga_on_failure,            --                   .boot_from_fpga_on_failure
			uart0_cts                     => hps_uart0_cts,                                      --              uart0.cts
			uart0_dsr                     => hps_uart0_dsr,                                      --                   .dsr
			uart0_dcd                     => hps_uart0_dcd,                                      --                   .dcd
			uart0_ri                      => hps_uart0_ri,                                       --                   .ri
			uart0_dtr                     => hps_uart0_dtr,                                      --                   .dtr
			uart0_rts                     => hps_uart0_rts,                                      --                   .rts
			uart0_out1_n                  => hps_uart0_out1_n,                                   --                   .out1_n
			uart0_out2_n                  => hps_uart0_out2_n,                                   --                   .out2_n
			uart0_rxd                     => hps_uart0_rxd,                                      --                   .rxd
			uart0_txd                     => hps_uart0_txd,                                      --                   .txd
			mem_a                         => memory_mem_a,                                       --             memory.mem_a
			mem_ba                        => memory_mem_ba,                                      --                   .mem_ba
			mem_ck                        => memory_mem_ck,                                      --                   .mem_ck
			mem_ck_n                      => memory_mem_ck_n,                                    --                   .mem_ck_n
			mem_cke                       => memory_mem_cke,                                     --                   .mem_cke
			mem_cs_n                      => memory_mem_cs_n,                                    --                   .mem_cs_n
			mem_ras_n                     => memory_mem_ras_n,                                   --                   .mem_ras_n
			mem_cas_n                     => memory_mem_cas_n,                                   --                   .mem_cas_n
			mem_we_n                      => memory_mem_we_n,                                    --                   .mem_we_n
			mem_reset_n                   => memory_mem_reset_n,                                 --                   .mem_reset_n
			mem_dq                        => memory_mem_dq,                                      --                   .mem_dq
			mem_dqs                       => memory_mem_dqs,                                     --                   .mem_dqs
			mem_dqs_n                     => memory_mem_dqs_n,                                   --                   .mem_dqs_n
			mem_odt                       => memory_mem_odt,                                     --                   .mem_odt
			mem_dm                        => memory_mem_dm,                                      --                   .mem_dm
			oct_rzqin                     => memory_oct_rzqin,                                   --                   .oct_rzqin
			hps_io_emac1_inst_TX_CLK      => hps_io_hps_io_emac1_inst_TX_CLK,                    --             hps_io.hps_io_emac1_inst_TX_CLK
			hps_io_emac1_inst_TXD0        => hps_io_hps_io_emac1_inst_TXD0,                      --                   .hps_io_emac1_inst_TXD0
			hps_io_emac1_inst_TXD1        => hps_io_hps_io_emac1_inst_TXD1,                      --                   .hps_io_emac1_inst_TXD1
			hps_io_emac1_inst_TXD2        => hps_io_hps_io_emac1_inst_TXD2,                      --                   .hps_io_emac1_inst_TXD2
			hps_io_emac1_inst_TXD3        => hps_io_hps_io_emac1_inst_TXD3,                      --                   .hps_io_emac1_inst_TXD3
			hps_io_emac1_inst_RXD0        => hps_io_hps_io_emac1_inst_RXD0,                      --                   .hps_io_emac1_inst_RXD0
			hps_io_emac1_inst_MDIO        => hps_io_hps_io_emac1_inst_MDIO,                      --                   .hps_io_emac1_inst_MDIO
			hps_io_emac1_inst_MDC         => hps_io_hps_io_emac1_inst_MDC,                       --                   .hps_io_emac1_inst_MDC
			hps_io_emac1_inst_RX_CTL      => hps_io_hps_io_emac1_inst_RX_CTL,                    --                   .hps_io_emac1_inst_RX_CTL
			hps_io_emac1_inst_TX_CTL      => hps_io_hps_io_emac1_inst_TX_CTL,                    --                   .hps_io_emac1_inst_TX_CTL
			hps_io_emac1_inst_RX_CLK      => hps_io_hps_io_emac1_inst_RX_CLK,                    --                   .hps_io_emac1_inst_RX_CLK
			hps_io_emac1_inst_RXD1        => hps_io_hps_io_emac1_inst_RXD1,                      --                   .hps_io_emac1_inst_RXD1
			hps_io_emac1_inst_RXD2        => hps_io_hps_io_emac1_inst_RXD2,                      --                   .hps_io_emac1_inst_RXD2
			hps_io_emac1_inst_RXD3        => hps_io_hps_io_emac1_inst_RXD3,                      --                   .hps_io_emac1_inst_RXD3
			hps_io_qspi_inst_IO0          => hps_io_hps_io_qspi_inst_IO0,                        --                   .hps_io_qspi_inst_IO0
			hps_io_qspi_inst_IO1          => hps_io_hps_io_qspi_inst_IO1,                        --                   .hps_io_qspi_inst_IO1
			hps_io_qspi_inst_IO2          => hps_io_hps_io_qspi_inst_IO2,                        --                   .hps_io_qspi_inst_IO2
			hps_io_qspi_inst_IO3          => hps_io_hps_io_qspi_inst_IO3,                        --                   .hps_io_qspi_inst_IO3
			hps_io_qspi_inst_SS0          => hps_io_hps_io_qspi_inst_SS0,                        --                   .hps_io_qspi_inst_SS0
			hps_io_qspi_inst_CLK          => hps_io_hps_io_qspi_inst_CLK,                        --                   .hps_io_qspi_inst_CLK
			hps_io_sdio_inst_CMD          => hps_io_hps_io_sdio_inst_CMD,                        --                   .hps_io_sdio_inst_CMD
			hps_io_sdio_inst_D0           => hps_io_hps_io_sdio_inst_D0,                         --                   .hps_io_sdio_inst_D0
			hps_io_sdio_inst_D1           => hps_io_hps_io_sdio_inst_D1,                         --                   .hps_io_sdio_inst_D1
			hps_io_sdio_inst_CLK          => hps_io_hps_io_sdio_inst_CLK,                        --                   .hps_io_sdio_inst_CLK
			hps_io_sdio_inst_D2           => hps_io_hps_io_sdio_inst_D2,                         --                   .hps_io_sdio_inst_D2
			hps_io_sdio_inst_D3           => hps_io_hps_io_sdio_inst_D3,                         --                   .hps_io_sdio_inst_D3
			hps_io_usb1_inst_D0           => hps_io_hps_io_usb1_inst_D0,                         --                   .hps_io_usb1_inst_D0
			hps_io_usb1_inst_D1           => hps_io_hps_io_usb1_inst_D1,                         --                   .hps_io_usb1_inst_D1
			hps_io_usb1_inst_D2           => hps_io_hps_io_usb1_inst_D2,                         --                   .hps_io_usb1_inst_D2
			hps_io_usb1_inst_D3           => hps_io_hps_io_usb1_inst_D3,                         --                   .hps_io_usb1_inst_D3
			hps_io_usb1_inst_D4           => hps_io_hps_io_usb1_inst_D4,                         --                   .hps_io_usb1_inst_D4
			hps_io_usb1_inst_D5           => hps_io_hps_io_usb1_inst_D5,                         --                   .hps_io_usb1_inst_D5
			hps_io_usb1_inst_D6           => hps_io_hps_io_usb1_inst_D6,                         --                   .hps_io_usb1_inst_D6
			hps_io_usb1_inst_D7           => hps_io_hps_io_usb1_inst_D7,                         --                   .hps_io_usb1_inst_D7
			hps_io_usb1_inst_CLK          => hps_io_hps_io_usb1_inst_CLK,                        --                   .hps_io_usb1_inst_CLK
			hps_io_usb1_inst_STP          => hps_io_hps_io_usb1_inst_STP,                        --                   .hps_io_usb1_inst_STP
			hps_io_usb1_inst_DIR          => hps_io_hps_io_usb1_inst_DIR,                        --                   .hps_io_usb1_inst_DIR
			hps_io_usb1_inst_NXT          => hps_io_hps_io_usb1_inst_NXT,                        --                   .hps_io_usb1_inst_NXT
			hps_io_spim1_inst_CLK         => hps_io_hps_io_spim1_inst_CLK,                       --                   .hps_io_spim1_inst_CLK
			hps_io_spim1_inst_MOSI        => hps_io_hps_io_spim1_inst_MOSI,                      --                   .hps_io_spim1_inst_MOSI
			hps_io_spim1_inst_MISO        => hps_io_hps_io_spim1_inst_MISO,                      --                   .hps_io_spim1_inst_MISO
			hps_io_spim1_inst_SS0         => hps_io_hps_io_spim1_inst_SS0,                       --                   .hps_io_spim1_inst_SS0
			hps_io_i2c0_inst_SDA          => hps_io_hps_io_i2c0_inst_SDA,                        --                   .hps_io_i2c0_inst_SDA
			hps_io_i2c0_inst_SCL          => hps_io_hps_io_i2c0_inst_SCL,                        --                   .hps_io_i2c0_inst_SCL
			hps_io_i2c1_inst_SDA          => hps_io_hps_io_i2c1_inst_SDA,                        --                   .hps_io_i2c1_inst_SDA
			hps_io_i2c1_inst_SCL          => hps_io_hps_io_i2c1_inst_SCL,                        --                   .hps_io_i2c1_inst_SCL
			hps_io_gpio_inst_GPIO09       => hps_io_hps_io_gpio_inst_GPIO09,                     --                   .hps_io_gpio_inst_GPIO09
			hps_io_gpio_inst_GPIO35       => hps_io_hps_io_gpio_inst_GPIO35,                     --                   .hps_io_gpio_inst_GPIO35
			hps_io_gpio_inst_GPIO40       => hps_io_hps_io_gpio_inst_GPIO40,                     --                   .hps_io_gpio_inst_GPIO40
			hps_io_gpio_inst_GPIO48       => hps_io_hps_io_gpio_inst_GPIO48,                     --                   .hps_io_gpio_inst_GPIO48
			hps_io_gpio_inst_GPIO61       => hps_io_hps_io_gpio_inst_GPIO61,                     --                   .hps_io_gpio_inst_GPIO61
			hps_io_gpio_inst_LOANIO49     => hps_io_hps_io_gpio_inst_LOANIO49,                   --                   .hps_io_gpio_inst_LOANIO49
			hps_io_gpio_inst_LOANIO50     => hps_io_hps_io_gpio_inst_LOANIO50,                   --                   .hps_io_gpio_inst_LOANIO50
			hps_io_gpio_inst_LOANIO53     => hps_io_hps_io_gpio_inst_LOANIO53,                   --                   .hps_io_gpio_inst_LOANIO53
			hps_io_gpio_inst_LOANIO54     => hps_io_hps_io_gpio_inst_LOANIO54,                   --                   .hps_io_gpio_inst_LOANIO54
			h2f_rst_n                     => arm_a9_hps_h2f_reset_reset,                         --          h2f_reset.reset_n
			h2f_axi_clk                   => system_pll_sys_clk_clk,                             --      h2f_axi_clock.clk
			h2f_AWID                      => arm_a9_hps_h2f_axi_master_awid,                     --     h2f_axi_master.awid
			h2f_AWADDR                    => arm_a9_hps_h2f_axi_master_awaddr,                   --                   .awaddr
			h2f_AWLEN                     => arm_a9_hps_h2f_axi_master_awlen,                    --                   .awlen
			h2f_AWSIZE                    => arm_a9_hps_h2f_axi_master_awsize,                   --                   .awsize
			h2f_AWBURST                   => arm_a9_hps_h2f_axi_master_awburst,                  --                   .awburst
			h2f_AWLOCK                    => arm_a9_hps_h2f_axi_master_awlock,                   --                   .awlock
			h2f_AWCACHE                   => arm_a9_hps_h2f_axi_master_awcache,                  --                   .awcache
			h2f_AWPROT                    => arm_a9_hps_h2f_axi_master_awprot,                   --                   .awprot
			h2f_AWVALID                   => arm_a9_hps_h2f_axi_master_awvalid,                  --                   .awvalid
			h2f_AWREADY                   => arm_a9_hps_h2f_axi_master_awready,                  --                   .awready
			h2f_WID                       => arm_a9_hps_h2f_axi_master_wid,                      --                   .wid
			h2f_WDATA                     => arm_a9_hps_h2f_axi_master_wdata,                    --                   .wdata
			h2f_WSTRB                     => arm_a9_hps_h2f_axi_master_wstrb,                    --                   .wstrb
			h2f_WLAST                     => arm_a9_hps_h2f_axi_master_wlast,                    --                   .wlast
			h2f_WVALID                    => arm_a9_hps_h2f_axi_master_wvalid,                   --                   .wvalid
			h2f_WREADY                    => arm_a9_hps_h2f_axi_master_wready,                   --                   .wready
			h2f_BID                       => arm_a9_hps_h2f_axi_master_bid,                      --                   .bid
			h2f_BRESP                     => arm_a9_hps_h2f_axi_master_bresp,                    --                   .bresp
			h2f_BVALID                    => arm_a9_hps_h2f_axi_master_bvalid,                   --                   .bvalid
			h2f_BREADY                    => arm_a9_hps_h2f_axi_master_bready,                   --                   .bready
			h2f_ARID                      => arm_a9_hps_h2f_axi_master_arid,                     --                   .arid
			h2f_ARADDR                    => arm_a9_hps_h2f_axi_master_araddr,                   --                   .araddr
			h2f_ARLEN                     => arm_a9_hps_h2f_axi_master_arlen,                    --                   .arlen
			h2f_ARSIZE                    => arm_a9_hps_h2f_axi_master_arsize,                   --                   .arsize
			h2f_ARBURST                   => arm_a9_hps_h2f_axi_master_arburst,                  --                   .arburst
			h2f_ARLOCK                    => arm_a9_hps_h2f_axi_master_arlock,                   --                   .arlock
			h2f_ARCACHE                   => arm_a9_hps_h2f_axi_master_arcache,                  --                   .arcache
			h2f_ARPROT                    => arm_a9_hps_h2f_axi_master_arprot,                   --                   .arprot
			h2f_ARVALID                   => arm_a9_hps_h2f_axi_master_arvalid,                  --                   .arvalid
			h2f_ARREADY                   => arm_a9_hps_h2f_axi_master_arready,                  --                   .arready
			h2f_RID                       => arm_a9_hps_h2f_axi_master_rid,                      --                   .rid
			h2f_RDATA                     => arm_a9_hps_h2f_axi_master_rdata,                    --                   .rdata
			h2f_RRESP                     => arm_a9_hps_h2f_axi_master_rresp,                    --                   .rresp
			h2f_RLAST                     => arm_a9_hps_h2f_axi_master_rlast,                    --                   .rlast
			h2f_RVALID                    => arm_a9_hps_h2f_axi_master_rvalid,                   --                   .rvalid
			h2f_RREADY                    => arm_a9_hps_h2f_axi_master_rready,                   --                   .rready
			f2h_axi_clk                   => system_pll_sys_clk_clk,                             --      f2h_axi_clock.clk
			f2h_AWID                      => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awid,    --      f2h_axi_slave.awid
			f2h_AWADDR                    => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awaddr,  --                   .awaddr
			f2h_AWLEN                     => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awlen,   --                   .awlen
			f2h_AWSIZE                    => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awsize,  --                   .awsize
			f2h_AWBURST                   => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awburst, --                   .awburst
			f2h_AWLOCK                    => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awlock,  --                   .awlock
			f2h_AWCACHE                   => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awcache, --                   .awcache
			f2h_AWPROT                    => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awprot,  --                   .awprot
			f2h_AWVALID                   => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awvalid, --                   .awvalid
			f2h_AWREADY                   => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awready, --                   .awready
			f2h_AWUSER                    => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awuser,  --                   .awuser
			f2h_WID                       => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wid,     --                   .wid
			f2h_WDATA                     => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wdata,   --                   .wdata
			f2h_WSTRB                     => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wstrb,   --                   .wstrb
			f2h_WLAST                     => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wlast,   --                   .wlast
			f2h_WVALID                    => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wvalid,  --                   .wvalid
			f2h_WREADY                    => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wready,  --                   .wready
			f2h_BID                       => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_bid,     --                   .bid
			f2h_BRESP                     => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_bresp,   --                   .bresp
			f2h_BVALID                    => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_bvalid,  --                   .bvalid
			f2h_BREADY                    => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_bready,  --                   .bready
			f2h_ARID                      => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arid,    --                   .arid
			f2h_ARADDR                    => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_araddr,  --                   .araddr
			f2h_ARLEN                     => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arlen,   --                   .arlen
			f2h_ARSIZE                    => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arsize,  --                   .arsize
			f2h_ARBURST                   => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arburst, --                   .arburst
			f2h_ARLOCK                    => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arlock,  --                   .arlock
			f2h_ARCACHE                   => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arcache, --                   .arcache
			f2h_ARPROT                    => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arprot,  --                   .arprot
			f2h_ARVALID                   => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arvalid, --                   .arvalid
			f2h_ARREADY                   => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arready, --                   .arready
			f2h_ARUSER                    => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_aruser,  --                   .aruser
			f2h_RID                       => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rid,     --                   .rid
			f2h_RDATA                     => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rdata,   --                   .rdata
			f2h_RRESP                     => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rresp,   --                   .rresp
			f2h_RLAST                     => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rlast,   --                   .rlast
			f2h_RVALID                    => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rvalid,  --                   .rvalid
			f2h_RREADY                    => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rready,  --                   .rready
			h2f_lw_axi_clk                => system_pll_sys_clk_clk,                             --   h2f_lw_axi_clock.clk
			h2f_lw_AWID                   => arm_a9_hps_h2f_lw_axi_master_awid,                  --  h2f_lw_axi_master.awid
			h2f_lw_AWADDR                 => arm_a9_hps_h2f_lw_axi_master_awaddr,                --                   .awaddr
			h2f_lw_AWLEN                  => arm_a9_hps_h2f_lw_axi_master_awlen,                 --                   .awlen
			h2f_lw_AWSIZE                 => arm_a9_hps_h2f_lw_axi_master_awsize,                --                   .awsize
			h2f_lw_AWBURST                => arm_a9_hps_h2f_lw_axi_master_awburst,               --                   .awburst
			h2f_lw_AWLOCK                 => arm_a9_hps_h2f_lw_axi_master_awlock,                --                   .awlock
			h2f_lw_AWCACHE                => arm_a9_hps_h2f_lw_axi_master_awcache,               --                   .awcache
			h2f_lw_AWPROT                 => arm_a9_hps_h2f_lw_axi_master_awprot,                --                   .awprot
			h2f_lw_AWVALID                => arm_a9_hps_h2f_lw_axi_master_awvalid,               --                   .awvalid
			h2f_lw_AWREADY                => arm_a9_hps_h2f_lw_axi_master_awready,               --                   .awready
			h2f_lw_WID                    => arm_a9_hps_h2f_lw_axi_master_wid,                   --                   .wid
			h2f_lw_WDATA                  => arm_a9_hps_h2f_lw_axi_master_wdata,                 --                   .wdata
			h2f_lw_WSTRB                  => arm_a9_hps_h2f_lw_axi_master_wstrb,                 --                   .wstrb
			h2f_lw_WLAST                  => arm_a9_hps_h2f_lw_axi_master_wlast,                 --                   .wlast
			h2f_lw_WVALID                 => arm_a9_hps_h2f_lw_axi_master_wvalid,                --                   .wvalid
			h2f_lw_WREADY                 => arm_a9_hps_h2f_lw_axi_master_wready,                --                   .wready
			h2f_lw_BID                    => arm_a9_hps_h2f_lw_axi_master_bid,                   --                   .bid
			h2f_lw_BRESP                  => arm_a9_hps_h2f_lw_axi_master_bresp,                 --                   .bresp
			h2f_lw_BVALID                 => arm_a9_hps_h2f_lw_axi_master_bvalid,                --                   .bvalid
			h2f_lw_BREADY                 => arm_a9_hps_h2f_lw_axi_master_bready,                --                   .bready
			h2f_lw_ARID                   => arm_a9_hps_h2f_lw_axi_master_arid,                  --                   .arid
			h2f_lw_ARADDR                 => arm_a9_hps_h2f_lw_axi_master_araddr,                --                   .araddr
			h2f_lw_ARLEN                  => arm_a9_hps_h2f_lw_axi_master_arlen,                 --                   .arlen
			h2f_lw_ARSIZE                 => arm_a9_hps_h2f_lw_axi_master_arsize,                --                   .arsize
			h2f_lw_ARBURST                => arm_a9_hps_h2f_lw_axi_master_arburst,               --                   .arburst
			h2f_lw_ARLOCK                 => arm_a9_hps_h2f_lw_axi_master_arlock,                --                   .arlock
			h2f_lw_ARCACHE                => arm_a9_hps_h2f_lw_axi_master_arcache,               --                   .arcache
			h2f_lw_ARPROT                 => arm_a9_hps_h2f_lw_axi_master_arprot,                --                   .arprot
			h2f_lw_ARVALID                => arm_a9_hps_h2f_lw_axi_master_arvalid,               --                   .arvalid
			h2f_lw_ARREADY                => arm_a9_hps_h2f_lw_axi_master_arready,               --                   .arready
			h2f_lw_RID                    => arm_a9_hps_h2f_lw_axi_master_rid,                   --                   .rid
			h2f_lw_RDATA                  => arm_a9_hps_h2f_lw_axi_master_rdata,                 --                   .rdata
			h2f_lw_RRESP                  => arm_a9_hps_h2f_lw_axi_master_rresp,                 --                   .rresp
			h2f_lw_RLAST                  => arm_a9_hps_h2f_lw_axi_master_rlast,                 --                   .rlast
			h2f_lw_RVALID                 => arm_a9_hps_h2f_lw_axi_master_rvalid,                --                   .rvalid
			h2f_lw_RREADY                 => arm_a9_hps_h2f_lw_axi_master_rready,                --                   .rready
			f2h_irq_p0                    => arm_a9_hps_f2h_irq0_irq,                            --           f2h_irq0.irq
			f2h_irq_p1                    => arm_a9_hps_f2h_irq1_irq                             --           f2h_irq1.irq
		);

	fpga_boot_sram : component Computer_System_FPGA_Boot_SRAM
		port map (
			clk        => system_pll_sys_clk_clk,                         --   clk1.clk
			address    => mm_interconnect_0_fpga_boot_sram_s1_address,    --     s1.address
			clken      => mm_interconnect_0_fpga_boot_sram_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_fpga_boot_sram_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_fpga_boot_sram_s1_write,      --       .write
			readdata   => mm_interconnect_0_fpga_boot_sram_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_fpga_boot_sram_s1_writedata,  --       .writedata
			reset      => rst_controller_reset_out_reset,                 -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req              --       .reset_req
		);

	jtag_uart_for_arm_0 : component Computer_System_JTAG_UART_for_ARM_0
		port map (
			clk            => system_pll_sys_clk_clk,                                                  --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                                --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_for_arm_0_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_for_arm_0_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_for_arm_0_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_for_arm_0_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_for_arm_0_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_for_arm_0_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_for_arm_0_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                                 --               irq.irq
		);

	jtag_uart_for_arm_1 : component Computer_System_JTAG_UART_for_ARM_0
		port map (
			clk            => system_pll_sys_clk_clk,                                                  --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                                --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_for_arm_1_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_for_arm_1_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_for_arm_1_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_for_arm_1_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_for_arm_1_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_for_arm_1_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_for_arm_1_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_001_receiver0_irq                                             --               irq.irq
		);

	jtag_to_fpga_bridge : component Computer_System_JTAG_to_FPGA_Bridge
		generic map (
			USE_PLI     => 0,
			PLI_PORT    => 50000,
			FIFO_DEPTHS => 2
		)
		port map (
			clk_clk              => system_pll_sys_clk_clk,                   --          clk.clk
			clk_reset_reset      => system_pll_reset_source_reset,            --    clk_reset.reset
			master_address       => jtag_to_fpga_bridge_master_address,       --       master.address
			master_readdata      => jtag_to_fpga_bridge_master_readdata,      --             .readdata
			master_read          => jtag_to_fpga_bridge_master_read,          --             .read
			master_write         => jtag_to_fpga_bridge_master_write,         --             .write
			master_writedata     => jtag_to_fpga_bridge_master_writedata,     --             .writedata
			master_waitrequest   => jtag_to_fpga_bridge_master_waitrequest,   --             .waitrequest
			master_readdatavalid => jtag_to_fpga_bridge_master_readdatavalid, --             .readdatavalid
			master_byteenable    => jtag_to_fpga_bridge_master_byteenable,    --             .byteenable
			master_reset_reset   => open                                      -- master_reset.reset
		);

	jtag_to_hps_bridge : component Computer_System_JTAG_to_FPGA_Bridge
		generic map (
			USE_PLI     => 0,
			PLI_PORT    => 50000,
			FIFO_DEPTHS => 2
		)
		port map (
			clk_clk              => system_pll_sys_clk_clk,                  --          clk.clk
			clk_reset_reset      => system_pll_reset_source_reset,           --    clk_reset.reset
			master_address       => jtag_to_hps_bridge_master_address,       --       master.address
			master_readdata      => jtag_to_hps_bridge_master_readdata,      --             .readdata
			master_read          => jtag_to_hps_bridge_master_read,          --             .read
			master_write         => jtag_to_hps_bridge_master_write,         --             .write
			master_writedata     => jtag_to_hps_bridge_master_writedata,     --             .writedata
			master_waitrequest   => jtag_to_hps_bridge_master_waitrequest,   --             .waitrequest
			master_readdatavalid => jtag_to_hps_bridge_master_readdatavalid, --             .readdatavalid
			master_byteenable    => jtag_to_hps_bridge_master_byteenable,    --             .byteenable
			master_reset_reset   => open                                     -- master_reset.reset
		);

	sysid : component Computer_System_SysID
		port map (
			clock    => system_pll_sys_clk_clk,                           --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,         --         reset.reset_n
			readdata => mm_interconnect_0_sysid_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_control_slave_address(0)  --              .address
		);

	system_pll : component Computer_System_System_PLL
		port map (
			ref_clk_clk        => system_clk_clk,                --      ref_clk.clk
			ref_reset_reset    => system_reset_reset,            --    ref_reset.reset
			sys_clk_clk        => system_pll_sys_clk_clk,        --      sys_clk.clk
			sdram_clk_clk      => open,                          --    sdram_clk.clk
			reset_source_reset => system_pll_reset_source_reset  -- reset_source.reset
		);

	mm_interconnect_0 : component Computer_System_mm_interconnect_0
		port map (
			ARM_A9_HPS_h2f_axi_master_awid                                        => arm_a9_hps_h2f_axi_master_awid,                                      --                                       ARM_A9_HPS_h2f_axi_master.awid
			ARM_A9_HPS_h2f_axi_master_awaddr                                      => arm_a9_hps_h2f_axi_master_awaddr,                                    --                                                                .awaddr
			ARM_A9_HPS_h2f_axi_master_awlen                                       => arm_a9_hps_h2f_axi_master_awlen,                                     --                                                                .awlen
			ARM_A9_HPS_h2f_axi_master_awsize                                      => arm_a9_hps_h2f_axi_master_awsize,                                    --                                                                .awsize
			ARM_A9_HPS_h2f_axi_master_awburst                                     => arm_a9_hps_h2f_axi_master_awburst,                                   --                                                                .awburst
			ARM_A9_HPS_h2f_axi_master_awlock                                      => arm_a9_hps_h2f_axi_master_awlock,                                    --                                                                .awlock
			ARM_A9_HPS_h2f_axi_master_awcache                                     => arm_a9_hps_h2f_axi_master_awcache,                                   --                                                                .awcache
			ARM_A9_HPS_h2f_axi_master_awprot                                      => arm_a9_hps_h2f_axi_master_awprot,                                    --                                                                .awprot
			ARM_A9_HPS_h2f_axi_master_awvalid                                     => arm_a9_hps_h2f_axi_master_awvalid,                                   --                                                                .awvalid
			ARM_A9_HPS_h2f_axi_master_awready                                     => arm_a9_hps_h2f_axi_master_awready,                                   --                                                                .awready
			ARM_A9_HPS_h2f_axi_master_wid                                         => arm_a9_hps_h2f_axi_master_wid,                                       --                                                                .wid
			ARM_A9_HPS_h2f_axi_master_wdata                                       => arm_a9_hps_h2f_axi_master_wdata,                                     --                                                                .wdata
			ARM_A9_HPS_h2f_axi_master_wstrb                                       => arm_a9_hps_h2f_axi_master_wstrb,                                     --                                                                .wstrb
			ARM_A9_HPS_h2f_axi_master_wlast                                       => arm_a9_hps_h2f_axi_master_wlast,                                     --                                                                .wlast
			ARM_A9_HPS_h2f_axi_master_wvalid                                      => arm_a9_hps_h2f_axi_master_wvalid,                                    --                                                                .wvalid
			ARM_A9_HPS_h2f_axi_master_wready                                      => arm_a9_hps_h2f_axi_master_wready,                                    --                                                                .wready
			ARM_A9_HPS_h2f_axi_master_bid                                         => arm_a9_hps_h2f_axi_master_bid,                                       --                                                                .bid
			ARM_A9_HPS_h2f_axi_master_bresp                                       => arm_a9_hps_h2f_axi_master_bresp,                                     --                                                                .bresp
			ARM_A9_HPS_h2f_axi_master_bvalid                                      => arm_a9_hps_h2f_axi_master_bvalid,                                    --                                                                .bvalid
			ARM_A9_HPS_h2f_axi_master_bready                                      => arm_a9_hps_h2f_axi_master_bready,                                    --                                                                .bready
			ARM_A9_HPS_h2f_axi_master_arid                                        => arm_a9_hps_h2f_axi_master_arid,                                      --                                                                .arid
			ARM_A9_HPS_h2f_axi_master_araddr                                      => arm_a9_hps_h2f_axi_master_araddr,                                    --                                                                .araddr
			ARM_A9_HPS_h2f_axi_master_arlen                                       => arm_a9_hps_h2f_axi_master_arlen,                                     --                                                                .arlen
			ARM_A9_HPS_h2f_axi_master_arsize                                      => arm_a9_hps_h2f_axi_master_arsize,                                    --                                                                .arsize
			ARM_A9_HPS_h2f_axi_master_arburst                                     => arm_a9_hps_h2f_axi_master_arburst,                                   --                                                                .arburst
			ARM_A9_HPS_h2f_axi_master_arlock                                      => arm_a9_hps_h2f_axi_master_arlock,                                    --                                                                .arlock
			ARM_A9_HPS_h2f_axi_master_arcache                                     => arm_a9_hps_h2f_axi_master_arcache,                                   --                                                                .arcache
			ARM_A9_HPS_h2f_axi_master_arprot                                      => arm_a9_hps_h2f_axi_master_arprot,                                    --                                                                .arprot
			ARM_A9_HPS_h2f_axi_master_arvalid                                     => arm_a9_hps_h2f_axi_master_arvalid,                                   --                                                                .arvalid
			ARM_A9_HPS_h2f_axi_master_arready                                     => arm_a9_hps_h2f_axi_master_arready,                                   --                                                                .arready
			ARM_A9_HPS_h2f_axi_master_rid                                         => arm_a9_hps_h2f_axi_master_rid,                                       --                                                                .rid
			ARM_A9_HPS_h2f_axi_master_rdata                                       => arm_a9_hps_h2f_axi_master_rdata,                                     --                                                                .rdata
			ARM_A9_HPS_h2f_axi_master_rresp                                       => arm_a9_hps_h2f_axi_master_rresp,                                     --                                                                .rresp
			ARM_A9_HPS_h2f_axi_master_rlast                                       => arm_a9_hps_h2f_axi_master_rlast,                                     --                                                                .rlast
			ARM_A9_HPS_h2f_axi_master_rvalid                                      => arm_a9_hps_h2f_axi_master_rvalid,                                    --                                                                .rvalid
			ARM_A9_HPS_h2f_axi_master_rready                                      => arm_a9_hps_h2f_axi_master_rready,                                    --                                                                .rready
			ARM_A9_HPS_h2f_lw_axi_master_awid                                     => arm_a9_hps_h2f_lw_axi_master_awid,                                   --                                    ARM_A9_HPS_h2f_lw_axi_master.awid
			ARM_A9_HPS_h2f_lw_axi_master_awaddr                                   => arm_a9_hps_h2f_lw_axi_master_awaddr,                                 --                                                                .awaddr
			ARM_A9_HPS_h2f_lw_axi_master_awlen                                    => arm_a9_hps_h2f_lw_axi_master_awlen,                                  --                                                                .awlen
			ARM_A9_HPS_h2f_lw_axi_master_awsize                                   => arm_a9_hps_h2f_lw_axi_master_awsize,                                 --                                                                .awsize
			ARM_A9_HPS_h2f_lw_axi_master_awburst                                  => arm_a9_hps_h2f_lw_axi_master_awburst,                                --                                                                .awburst
			ARM_A9_HPS_h2f_lw_axi_master_awlock                                   => arm_a9_hps_h2f_lw_axi_master_awlock,                                 --                                                                .awlock
			ARM_A9_HPS_h2f_lw_axi_master_awcache                                  => arm_a9_hps_h2f_lw_axi_master_awcache,                                --                                                                .awcache
			ARM_A9_HPS_h2f_lw_axi_master_awprot                                   => arm_a9_hps_h2f_lw_axi_master_awprot,                                 --                                                                .awprot
			ARM_A9_HPS_h2f_lw_axi_master_awvalid                                  => arm_a9_hps_h2f_lw_axi_master_awvalid,                                --                                                                .awvalid
			ARM_A9_HPS_h2f_lw_axi_master_awready                                  => arm_a9_hps_h2f_lw_axi_master_awready,                                --                                                                .awready
			ARM_A9_HPS_h2f_lw_axi_master_wid                                      => arm_a9_hps_h2f_lw_axi_master_wid,                                    --                                                                .wid
			ARM_A9_HPS_h2f_lw_axi_master_wdata                                    => arm_a9_hps_h2f_lw_axi_master_wdata,                                  --                                                                .wdata
			ARM_A9_HPS_h2f_lw_axi_master_wstrb                                    => arm_a9_hps_h2f_lw_axi_master_wstrb,                                  --                                                                .wstrb
			ARM_A9_HPS_h2f_lw_axi_master_wlast                                    => arm_a9_hps_h2f_lw_axi_master_wlast,                                  --                                                                .wlast
			ARM_A9_HPS_h2f_lw_axi_master_wvalid                                   => arm_a9_hps_h2f_lw_axi_master_wvalid,                                 --                                                                .wvalid
			ARM_A9_HPS_h2f_lw_axi_master_wready                                   => arm_a9_hps_h2f_lw_axi_master_wready,                                 --                                                                .wready
			ARM_A9_HPS_h2f_lw_axi_master_bid                                      => arm_a9_hps_h2f_lw_axi_master_bid,                                    --                                                                .bid
			ARM_A9_HPS_h2f_lw_axi_master_bresp                                    => arm_a9_hps_h2f_lw_axi_master_bresp,                                  --                                                                .bresp
			ARM_A9_HPS_h2f_lw_axi_master_bvalid                                   => arm_a9_hps_h2f_lw_axi_master_bvalid,                                 --                                                                .bvalid
			ARM_A9_HPS_h2f_lw_axi_master_bready                                   => arm_a9_hps_h2f_lw_axi_master_bready,                                 --                                                                .bready
			ARM_A9_HPS_h2f_lw_axi_master_arid                                     => arm_a9_hps_h2f_lw_axi_master_arid,                                   --                                                                .arid
			ARM_A9_HPS_h2f_lw_axi_master_araddr                                   => arm_a9_hps_h2f_lw_axi_master_araddr,                                 --                                                                .araddr
			ARM_A9_HPS_h2f_lw_axi_master_arlen                                    => arm_a9_hps_h2f_lw_axi_master_arlen,                                  --                                                                .arlen
			ARM_A9_HPS_h2f_lw_axi_master_arsize                                   => arm_a9_hps_h2f_lw_axi_master_arsize,                                 --                                                                .arsize
			ARM_A9_HPS_h2f_lw_axi_master_arburst                                  => arm_a9_hps_h2f_lw_axi_master_arburst,                                --                                                                .arburst
			ARM_A9_HPS_h2f_lw_axi_master_arlock                                   => arm_a9_hps_h2f_lw_axi_master_arlock,                                 --                                                                .arlock
			ARM_A9_HPS_h2f_lw_axi_master_arcache                                  => arm_a9_hps_h2f_lw_axi_master_arcache,                                --                                                                .arcache
			ARM_A9_HPS_h2f_lw_axi_master_arprot                                   => arm_a9_hps_h2f_lw_axi_master_arprot,                                 --                                                                .arprot
			ARM_A9_HPS_h2f_lw_axi_master_arvalid                                  => arm_a9_hps_h2f_lw_axi_master_arvalid,                                --                                                                .arvalid
			ARM_A9_HPS_h2f_lw_axi_master_arready                                  => arm_a9_hps_h2f_lw_axi_master_arready,                                --                                                                .arready
			ARM_A9_HPS_h2f_lw_axi_master_rid                                      => arm_a9_hps_h2f_lw_axi_master_rid,                                    --                                                                .rid
			ARM_A9_HPS_h2f_lw_axi_master_rdata                                    => arm_a9_hps_h2f_lw_axi_master_rdata,                                  --                                                                .rdata
			ARM_A9_HPS_h2f_lw_axi_master_rresp                                    => arm_a9_hps_h2f_lw_axi_master_rresp,                                  --                                                                .rresp
			ARM_A9_HPS_h2f_lw_axi_master_rlast                                    => arm_a9_hps_h2f_lw_axi_master_rlast,                                  --                                                                .rlast
			ARM_A9_HPS_h2f_lw_axi_master_rvalid                                   => arm_a9_hps_h2f_lw_axi_master_rvalid,                                 --                                                                .rvalid
			ARM_A9_HPS_h2f_lw_axi_master_rready                                   => arm_a9_hps_h2f_lw_axi_master_rready,                                 --                                                                .rready
			System_PLL_sys_clk_clk                                                => system_pll_sys_clk_clk,                                              --                                              System_PLL_sys_clk.clk
			ARM_A9_HPS_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,                                  -- ARM_A9_HPS_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
			FPGA_Boot_SRAM_reset1_reset_bridge_in_reset_reset                     => rst_controller_reset_out_reset,                                      --                     FPGA_Boot_SRAM_reset1_reset_bridge_in_reset.reset
			JTAG_to_FPGA_Bridge_clk_reset_reset_bridge_in_reset_reset             => rst_controller_reset_out_reset,                                      --             JTAG_to_FPGA_Bridge_clk_reset_reset_bridge_in_reset.reset
			JTAG_to_FPGA_Bridge_master_address                                    => jtag_to_fpga_bridge_master_address,                                  --                                      JTAG_to_FPGA_Bridge_master.address
			JTAG_to_FPGA_Bridge_master_waitrequest                                => jtag_to_fpga_bridge_master_waitrequest,                              --                                                                .waitrequest
			JTAG_to_FPGA_Bridge_master_byteenable                                 => jtag_to_fpga_bridge_master_byteenable,                               --                                                                .byteenable
			JTAG_to_FPGA_Bridge_master_read                                       => jtag_to_fpga_bridge_master_read,                                     --                                                                .read
			JTAG_to_FPGA_Bridge_master_readdata                                   => jtag_to_fpga_bridge_master_readdata,                                 --                                                                .readdata
			JTAG_to_FPGA_Bridge_master_readdatavalid                              => jtag_to_fpga_bridge_master_readdatavalid,                            --                                                                .readdatavalid
			JTAG_to_FPGA_Bridge_master_write                                      => jtag_to_fpga_bridge_master_write,                                    --                                                                .write
			JTAG_to_FPGA_Bridge_master_writedata                                  => jtag_to_fpga_bridge_master_writedata,                                --                                                                .writedata
			FPGA_Boot_SRAM_s1_address                                             => mm_interconnect_0_fpga_boot_sram_s1_address,                         --                                               FPGA_Boot_SRAM_s1.address
			FPGA_Boot_SRAM_s1_write                                               => mm_interconnect_0_fpga_boot_sram_s1_write,                           --                                                                .write
			FPGA_Boot_SRAM_s1_readdata                                            => mm_interconnect_0_fpga_boot_sram_s1_readdata,                        --                                                                .readdata
			FPGA_Boot_SRAM_s1_writedata                                           => mm_interconnect_0_fpga_boot_sram_s1_writedata,                       --                                                                .writedata
			FPGA_Boot_SRAM_s1_chipselect                                          => mm_interconnect_0_fpga_boot_sram_s1_chipselect,                      --                                                                .chipselect
			FPGA_Boot_SRAM_s1_clken                                               => mm_interconnect_0_fpga_boot_sram_s1_clken,                           --                                                                .clken
			JTAG_UART_for_ARM_0_avalon_jtag_slave_address                         => mm_interconnect_0_jtag_uart_for_arm_0_avalon_jtag_slave_address,     --                           JTAG_UART_for_ARM_0_avalon_jtag_slave.address
			JTAG_UART_for_ARM_0_avalon_jtag_slave_write                           => mm_interconnect_0_jtag_uart_for_arm_0_avalon_jtag_slave_write,       --                                                                .write
			JTAG_UART_for_ARM_0_avalon_jtag_slave_read                            => mm_interconnect_0_jtag_uart_for_arm_0_avalon_jtag_slave_read,        --                                                                .read
			JTAG_UART_for_ARM_0_avalon_jtag_slave_readdata                        => mm_interconnect_0_jtag_uart_for_arm_0_avalon_jtag_slave_readdata,    --                                                                .readdata
			JTAG_UART_for_ARM_0_avalon_jtag_slave_writedata                       => mm_interconnect_0_jtag_uart_for_arm_0_avalon_jtag_slave_writedata,   --                                                                .writedata
			JTAG_UART_for_ARM_0_avalon_jtag_slave_waitrequest                     => mm_interconnect_0_jtag_uart_for_arm_0_avalon_jtag_slave_waitrequest, --                                                                .waitrequest
			JTAG_UART_for_ARM_0_avalon_jtag_slave_chipselect                      => mm_interconnect_0_jtag_uart_for_arm_0_avalon_jtag_slave_chipselect,  --                                                                .chipselect
			JTAG_UART_for_ARM_1_avalon_jtag_slave_address                         => mm_interconnect_0_jtag_uart_for_arm_1_avalon_jtag_slave_address,     --                           JTAG_UART_for_ARM_1_avalon_jtag_slave.address
			JTAG_UART_for_ARM_1_avalon_jtag_slave_write                           => mm_interconnect_0_jtag_uart_for_arm_1_avalon_jtag_slave_write,       --                                                                .write
			JTAG_UART_for_ARM_1_avalon_jtag_slave_read                            => mm_interconnect_0_jtag_uart_for_arm_1_avalon_jtag_slave_read,        --                                                                .read
			JTAG_UART_for_ARM_1_avalon_jtag_slave_readdata                        => mm_interconnect_0_jtag_uart_for_arm_1_avalon_jtag_slave_readdata,    --                                                                .readdata
			JTAG_UART_for_ARM_1_avalon_jtag_slave_writedata                       => mm_interconnect_0_jtag_uart_for_arm_1_avalon_jtag_slave_writedata,   --                                                                .writedata
			JTAG_UART_for_ARM_1_avalon_jtag_slave_waitrequest                     => mm_interconnect_0_jtag_uart_for_arm_1_avalon_jtag_slave_waitrequest, --                                                                .waitrequest
			JTAG_UART_for_ARM_1_avalon_jtag_slave_chipselect                      => mm_interconnect_0_jtag_uart_for_arm_1_avalon_jtag_slave_chipselect,  --                                                                .chipselect
			SysID_control_slave_address                                           => mm_interconnect_0_sysid_control_slave_address,                       --                                             SysID_control_slave.address
			SysID_control_slave_readdata                                          => mm_interconnect_0_sysid_control_slave_readdata                       --                                                                .readdata
		);

	mm_interconnect_1 : component Computer_System_mm_interconnect_1
		port map (
			ARM_A9_HPS_f2h_axi_slave_awid                                          => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awid,    --                                         ARM_A9_HPS_f2h_axi_slave.awid
			ARM_A9_HPS_f2h_axi_slave_awaddr                                        => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awaddr,  --                                                                 .awaddr
			ARM_A9_HPS_f2h_axi_slave_awlen                                         => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awlen,   --                                                                 .awlen
			ARM_A9_HPS_f2h_axi_slave_awsize                                        => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awsize,  --                                                                 .awsize
			ARM_A9_HPS_f2h_axi_slave_awburst                                       => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awburst, --                                                                 .awburst
			ARM_A9_HPS_f2h_axi_slave_awlock                                        => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awlock,  --                                                                 .awlock
			ARM_A9_HPS_f2h_axi_slave_awcache                                       => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awcache, --                                                                 .awcache
			ARM_A9_HPS_f2h_axi_slave_awprot                                        => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awprot,  --                                                                 .awprot
			ARM_A9_HPS_f2h_axi_slave_awuser                                        => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awuser,  --                                                                 .awuser
			ARM_A9_HPS_f2h_axi_slave_awvalid                                       => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awvalid, --                                                                 .awvalid
			ARM_A9_HPS_f2h_axi_slave_awready                                       => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_awready, --                                                                 .awready
			ARM_A9_HPS_f2h_axi_slave_wid                                           => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wid,     --                                                                 .wid
			ARM_A9_HPS_f2h_axi_slave_wdata                                         => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wdata,   --                                                                 .wdata
			ARM_A9_HPS_f2h_axi_slave_wstrb                                         => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wstrb,   --                                                                 .wstrb
			ARM_A9_HPS_f2h_axi_slave_wlast                                         => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wlast,   --                                                                 .wlast
			ARM_A9_HPS_f2h_axi_slave_wvalid                                        => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wvalid,  --                                                                 .wvalid
			ARM_A9_HPS_f2h_axi_slave_wready                                        => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_wready,  --                                                                 .wready
			ARM_A9_HPS_f2h_axi_slave_bid                                           => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_bid,     --                                                                 .bid
			ARM_A9_HPS_f2h_axi_slave_bresp                                         => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_bresp,   --                                                                 .bresp
			ARM_A9_HPS_f2h_axi_slave_bvalid                                        => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_bvalid,  --                                                                 .bvalid
			ARM_A9_HPS_f2h_axi_slave_bready                                        => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_bready,  --                                                                 .bready
			ARM_A9_HPS_f2h_axi_slave_arid                                          => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arid,    --                                                                 .arid
			ARM_A9_HPS_f2h_axi_slave_araddr                                        => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_araddr,  --                                                                 .araddr
			ARM_A9_HPS_f2h_axi_slave_arlen                                         => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arlen,   --                                                                 .arlen
			ARM_A9_HPS_f2h_axi_slave_arsize                                        => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arsize,  --                                                                 .arsize
			ARM_A9_HPS_f2h_axi_slave_arburst                                       => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arburst, --                                                                 .arburst
			ARM_A9_HPS_f2h_axi_slave_arlock                                        => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arlock,  --                                                                 .arlock
			ARM_A9_HPS_f2h_axi_slave_arcache                                       => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arcache, --                                                                 .arcache
			ARM_A9_HPS_f2h_axi_slave_arprot                                        => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arprot,  --                                                                 .arprot
			ARM_A9_HPS_f2h_axi_slave_aruser                                        => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_aruser,  --                                                                 .aruser
			ARM_A9_HPS_f2h_axi_slave_arvalid                                       => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arvalid, --                                                                 .arvalid
			ARM_A9_HPS_f2h_axi_slave_arready                                       => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_arready, --                                                                 .arready
			ARM_A9_HPS_f2h_axi_slave_rid                                           => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rid,     --                                                                 .rid
			ARM_A9_HPS_f2h_axi_slave_rdata                                         => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rdata,   --                                                                 .rdata
			ARM_A9_HPS_f2h_axi_slave_rresp                                         => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rresp,   --                                                                 .rresp
			ARM_A9_HPS_f2h_axi_slave_rlast                                         => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rlast,   --                                                                 .rlast
			ARM_A9_HPS_f2h_axi_slave_rvalid                                        => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rvalid,  --                                                                 .rvalid
			ARM_A9_HPS_f2h_axi_slave_rready                                        => mm_interconnect_1_arm_a9_hps_f2h_axi_slave_rready,  --                                                                 .rready
			System_PLL_sys_clk_clk                                                 => system_pll_sys_clk_clk,                             --                                               System_PLL_sys_clk.clk
			ARM_A9_HPS_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset_reset  => rst_controller_001_reset_out_reset,                 --  ARM_A9_HPS_f2h_axi_slave_agent_reset_sink_reset_bridge_in_reset.reset
			JTAG_to_HPS_Bridge_clk_reset_reset_bridge_in_reset_reset               => rst_controller_reset_out_reset,                     --               JTAG_to_HPS_Bridge_clk_reset_reset_bridge_in_reset.reset
			JTAG_to_HPS_Bridge_master_translator_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                     -- JTAG_to_HPS_Bridge_master_translator_reset_reset_bridge_in_reset.reset
			JTAG_to_HPS_Bridge_master_address                                      => jtag_to_hps_bridge_master_address,                  --                                        JTAG_to_HPS_Bridge_master.address
			JTAG_to_HPS_Bridge_master_waitrequest                                  => jtag_to_hps_bridge_master_waitrequest,              --                                                                 .waitrequest
			JTAG_to_HPS_Bridge_master_byteenable                                   => jtag_to_hps_bridge_master_byteenable,               --                                                                 .byteenable
			JTAG_to_HPS_Bridge_master_read                                         => jtag_to_hps_bridge_master_read,                     --                                                                 .read
			JTAG_to_HPS_Bridge_master_readdata                                     => jtag_to_hps_bridge_master_readdata,                 --                                                                 .readdata
			JTAG_to_HPS_Bridge_master_readdatavalid                                => jtag_to_hps_bridge_master_readdatavalid,            --                                                                 .readdatavalid
			JTAG_to_HPS_Bridge_master_write                                        => jtag_to_hps_bridge_master_write,                    --                                                                 .write
			JTAG_to_HPS_Bridge_master_writedata                                    => jtag_to_hps_bridge_master_writedata                 --                                                                 .writedata
		);

	irq_mapper : component Computer_System_irq_mapper
		port map (
			clk           => open,                     --       clk.clk
			reset         => open,                     -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq, -- receiver0.irq
			sender_irq    => arm_a9_hps_f2h_irq0_irq   --    sender.irq
		);

	irq_mapper_001 : component Computer_System_irq_mapper
		port map (
			clk           => open,                         --       clk.clk
			reset         => open,                         -- clk_reset.reset
			receiver0_irq => irq_mapper_001_receiver0_irq, -- receiver0.irq
			sender_irq    => arm_a9_hps_f2h_irq1_irq       --    sender.irq
		);

	rst_controller : component computer_system_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => system_pll_reset_source_reset,      -- reset_in0.reset
			clk            => system_pll_sys_clk_clk,             --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_001 : component computer_system_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => fpga_reset_reset_n_ports_inv,       -- reset_in0.reset
			clk            => system_pll_sys_clk_clk,             --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	fpga_reset_reset_n_ports_inv <= not arm_a9_hps_h2f_reset_reset;

	mm_interconnect_0_jtag_uart_for_arm_0_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_for_arm_0_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_for_arm_0_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_for_arm_0_avalon_jtag_slave_write;

	mm_interconnect_0_jtag_uart_for_arm_1_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_for_arm_1_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_for_arm_1_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_for_arm_1_avalon_jtag_slave_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	fpga_reset_reset_n <= arm_a9_hps_h2f_reset_reset;

end architecture rtl; -- of Computer_System
