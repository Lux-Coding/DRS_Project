--------------------------------------------------------------------------------
-- Title       : HPS instantiation helper
-- Project     : FPGA Based Digital Signal Processing
--               FH OÖ Hagenberg/HSD, SCD5
--------------------------------------------------------------------------------
-- RevCtrl     : $Id: HPSComputerMin-e.vhd 733 2017-12-04 02:28:35Z mroland $
-- Authors     : Michael Roland, Hagenberg/Austria, Copyright (c) 2016-2017
--------------------------------------------------------------------------------
-- Description : Minimal Hard Prosessor System SoC Instantiation for access to
--               UART pins of HPS on Altera DE1-SoC
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.global.all;

entity HPSComputerMin is

  generic (
    gSimulationResetDeassertAfter : time := 117 ns
  );
  
  port (
    -- CLOCK
    CLOCK_50         : in    std_ulogic;
    
    -- RESET (for FPGA, generated by HPS)
    FPGA_RESET_N     : out   std_ulogic;
    
    -- UART (HPS LOAN I/O -> FPGA)
    FPGA_UART_TX     : in    std_ulogic;
    FPGA_UART_RX     : out   std_ulogic;
    
    -- HPS GPIO DEBUG
    MIRROR_HPS_LED   : out   std_ulogic;
    
    ----------------------------------------------------------------------------
    -- HPS I/O PINS
    ----------------------------------------------------------------------------
    
    -- DDR3 SDRAM
    HPS_DDR3_ADDR    : out   std_logic_vector(14 downto 0);
    HPS_DDR3_BA      : out   std_logic_vector(2 downto 0);
    HPS_DDR3_CK_P    : out   std_logic;
    HPS_DDR3_CK_N    : out   std_logic;
    HPS_DDR3_CKE     : out   std_logic;
    HPS_DDR3_CS_N    : out   std_logic;
    HPS_DDR3_RAS_N   : out   std_logic;
    HPS_DDR3_CAS_N   : out   std_logic;
    HPS_DDR3_WE_N    : out   std_logic;
    HPS_DDR3_RESET_N : out   std_logic;
    HPS_DDR3_DQ      : inout std_logic_vector(31 downto 0);
    HPS_DDR3_DQS_P   : inout std_logic_vector(3 downto 0);
    HPS_DDR3_DQS_N   : inout std_logic_vector(3 downto 0);
    HPS_DDR3_ODT     : out   std_logic;
    HPS_DDR3_DM      : out   std_logic_vector(3 downto 0);
    HPS_DDR3_RZQ     : in    std_logic;
    
    -- ETHERNET
    HPS_ENET_GTX_CLK : out   std_logic;
    HPS_ENET_MDC     : out   std_logic;
    HPS_ENET_MDIO    : inout std_logic;
    HPS_ENET_RX_CLK  : in    std_logic;
    HPS_ENET_RX_DATA : in    std_logic_vector(3 downto 0);
    HPS_ENET_RX_DV   : in    std_logic;
    HPS_ENET_TX_DATA : out   std_logic_vector(3 downto 0);
    HPS_ENET_TX_EN   : out   std_logic;
    HPS_ENET_INT_N   : inout std_logic;  -- HPS_GPIO35
    
    -- QSPI FLASH
    HPS_FLASH_DATA   : inout std_logic_vector(3 downto 0);
    HPS_FLASH_DCLK   : out   std_logic;
    HPS_FLASH_NCSO   : out   std_logic;
    
    -- I2C
    HPS_I2C_CONTROL  : inout std_logic;  -- HPS_GPIO48
    HPS_I2C1_SCLK    : inout std_logic;
    HPS_I2C1_SDAT    : inout std_logic;
    HPS_I2C2_SCLK    : inout std_logic;
    HPS_I2C2_SDAT    : inout std_logic;
    
    -- SD CARD
    HPS_SD_CMD       : inout std_logic;
    HPS_SD_CLK       : out   std_logic;
    HPS_SD_DATA      : inout std_logic_vector(3 downto 0);
    
    -- USB
    HPS_USB_CLKOUT   : in    std_logic;
    HPS_USB_DATA     : inout std_logic_vector(7 downto 0);
    HPS_USB_DIR      : in    std_logic;
    HPS_USB_NXT      : in    std_logic;
    HPS_USB_STP      : out   std_logic;
    HPS_CONV_USB_N   : inout std_logic;  -- HPS_GPIO09
    
    -- SPI
    HPS_SPIM_CLK     : out   std_logic;
    HPS_SPIM_MISO    : in    std_logic;
    HPS_SPIM_MOSI    : out   std_logic;
    HPS_SPIM_SS      : out   std_logic;

    -- UART
    HPS_UART_TX      : inout std_logic;  -- HPS_GPIO50
    HPS_UART_RX      : inout std_logic;  -- HPS_GPIO49
    
    -- GPIO
    HPS_KEY          : inout std_logic;  -- HPS_GPIO54
    HPS_LED          : inout std_logic;  -- HPS_GPIO53
    HPS_LTC_GPIO     : inout std_logic;  -- HPS_GPIO40
    HPS_GSENSOR_INT  : inout std_logic); -- HPS_GPIO61

end HPSComputerMin;
